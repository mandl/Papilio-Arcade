-- generated with romgen v3.04 by MikeJ
-- dummy rom. random rom data. avoid map to optimise this rom away;
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

--library UNISIM;
	--use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
port (
	CLK  : in  std_logic;
	ADDR : in  std_logic_vector(13 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_PGM_0 is


	type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
	signal ROM : ROM_ARRAY := (
		x"7A",x"B2",x"88",x"6A",x"94",x"C6",x"58",x"7F", -- 0x0000
		x"64",x"2E",x"AB",x"09",x"25",x"EB",x"52",x"C7", -- 0x0008
		x"0A",x"67",x"10",x"64",x"3A",x"B7",x"44",x"BA", -- 0x0010
		x"31",x"DB",x"63",x"30",x"6E",x"A4",x"80",x"69", -- 0x0018
		x"57",x"88",x"D3",x"6B",x"CF",x"2C",x"EA",x"B3", -- 0x0020
		x"D9",x"97",x"BC",x"FE",x"83",x"8F",x"47",x"0D", -- 0x0028
		x"76",x"D6",x"71",x"B0",x"8F",x"B5",x"EB",x"40", -- 0x0030
		x"12",x"4F",x"71",x"00",x"F3",x"F1",x"69",x"CA", -- 0x0038
		x"F9",x"BC",x"36",x"C9",x"68",x"22",x"FD",x"42", -- 0x0040
		x"39",x"3A",x"C1",x"3C",x"C9",x"09",x"49",x"41", -- 0x0048
		x"DF",x"3B",x"71",x"EE",x"70",x"5D",x"30",x"02", -- 0x0050
		x"AD",x"A1",x"03",x"21",x"13",x"EB",x"EC",x"0D", -- 0x0058
		x"A9",x"A2",x"57",x"91",x"C4",x"55",x"D4",x"7D", -- 0x0060
		x"8F",x"16",x"B9",x"5A",x"1F",x"83",x"1B",x"7E", -- 0x0068
		x"3E",x"8C",x"ED",x"AE",x"EA",x"1E",x"B1",x"18", -- 0x0070
		x"BF",x"34",x"39",x"D2",x"20",x"A5",x"5F",x"49", -- 0x0078
		x"49",x"B6",x"DB",x"8D",x"0C",x"30",x"0C",x"9C", -- 0x0080
		x"46",x"45",x"76",x"E4",x"48",x"91",x"E2",x"86", -- 0x0088
		x"9D",x"50",x"36",x"08",x"6E",x"67",x"20",x"AD", -- 0x0090
		x"9B",x"D9",x"80",x"3B",x"7F",x"E0",x"85",x"48", -- 0x0098
		x"97",x"E0",x"D6",x"24",x"90",x"62",x"40",x"56", -- 0x00A0
		x"27",x"B6",x"BA",x"70",x"C7",x"1D",x"76",x"E4", -- 0x00A8
		x"6E",x"2C",x"ED",x"DC",x"93",x"8D",x"8B",x"2F", -- 0x00B0
		x"67",x"8B",x"6B",x"67",x"EB",x"70",x"2F",x"04", -- 0x00B8
		x"D0",x"06",x"28",x"61",x"E7",x"68",x"B7",x"10", -- 0x00C0
		x"9E",x"F1",x"00",x"E5",x"0F",x"F5",x"CA",x"FC", -- 0x00C8
		x"23",x"B8",x"DA",x"B6",x"C6",x"E5",x"66",x"2E", -- 0x00D0
		x"F0",x"D1",x"15",x"DD",x"C1",x"45",x"E1",x"92", -- 0x00D8
		x"CA",x"89",x"F3",x"B3",x"F1",x"2B",x"43",x"10", -- 0x00E0
		x"1D",x"C2",x"F5",x"AB",x"B8",x"40",x"A9",x"5B", -- 0x00E8
		x"79",x"04",x"13",x"40",x"E9",x"79",x"ED",x"DA", -- 0x00F0
		x"CA",x"04",x"38",x"8C",x"C8",x"1A",x"1F",x"93", -- 0x00F8
		x"A3",x"92",x"C6",x"15",x"3D",x"89",x"25",x"D9", -- 0x0100
		x"CB",x"9A",x"85",x"05",x"DB",x"AE",x"60",x"55", -- 0x0108
		x"B2",x"73",x"15",x"1C",x"6C",x"03",x"77",x"37", -- 0x0110
		x"86",x"AF",x"43",x"4F",x"4A",x"E1",x"63",x"6D", -- 0x0118
		x"F3",x"A9",x"83",x"31",x"B3",x"28",x"0B",x"7F", -- 0x0120
		x"43",x"11",x"84",x"1F",x"BF",x"65",x"F3",x"F2", -- 0x0128
		x"58",x"09",x"0F",x"C5",x"0C",x"06",x"7C",x"13", -- 0x0130
		x"B6",x"40",x"62",x"80",x"22",x"45",x"ED",x"17", -- 0x0138
		x"EF",x"71",x"C7",x"A3",x"1A",x"D3",x"A2",x"5D", -- 0x0140
		x"E4",x"A7",x"FB",x"24",x"0D",x"EF",x"17",x"65", -- 0x0148
		x"78",x"A6",x"AA",x"04",x"AC",x"A7",x"17",x"E2", -- 0x0150
		x"E7",x"F9",x"63",x"89",x"3F",x"52",x"20",x"AE", -- 0x0158
		x"43",x"E8",x"52",x"5D",x"3C",x"F5",x"3A",x"A0", -- 0x0160
		x"1D",x"36",x"C4",x"2A",x"A5",x"DC",x"0F",x"1E", -- 0x0168
		x"83",x"BA",x"A2",x"AF",x"E1",x"B9",x"93",x"49", -- 0x0170
		x"33",x"F6",x"D2",x"73",x"C8",x"73",x"22",x"8C", -- 0x0178
		x"DB",x"F4",x"69",x"18",x"6A",x"A4",x"38",x"87", -- 0x0180
		x"5A",x"FC",x"31",x"01",x"59",x"40",x"9E",x"5C", -- 0x0188
		x"7A",x"41",x"0D",x"5C",x"7B",x"A0",x"A5",x"AE", -- 0x0190
		x"17",x"F8",x"A1",x"60",x"EB",x"44",x"EC",x"C7", -- 0x0198
		x"39",x"56",x"5F",x"23",x"7A",x"17",x"AA",x"D5", -- 0x01A0
		x"14",x"DB",x"56",x"ED",x"9B",x"74",x"4A",x"17", -- 0x01A8
		x"B6",x"D6",x"73",x"B1",x"F6",x"99",x"DF",x"8E", -- 0x01B0
		x"12",x"82",x"EE",x"FD",x"C6",x"5B",x"45",x"7F", -- 0x01B8
		x"31",x"24",x"A2",x"AC",x"3B",x"CC",x"02",x"CE", -- 0x01C0
		x"A8",x"D7",x"BC",x"44",x"4C",x"87",x"DA",x"82", -- 0x01C8
		x"5E",x"CE",x"34",x"56",x"68",x"15",x"E4",x"F9", -- 0x01D0
		x"17",x"53",x"77",x"DD",x"AE",x"BC",x"DC",x"DF", -- 0x01D8
		x"E0",x"FE",x"0C",x"9B",x"CB",x"8D",x"6A",x"74", -- 0x01E0
		x"65",x"A7",x"38",x"B2",x"2F",x"14",x"35",x"8D", -- 0x01E8
		x"E2",x"6A",x"63",x"CA",x"FE",x"C7",x"44",x"16", -- 0x01F0
		x"9A",x"BB",x"73",x"49",x"78",x"CF",x"A9",x"D8", -- 0x01F8
		x"CE",x"B5",x"74",x"9A",x"44",x"5E",x"8E",x"29", -- 0x0200
		x"06",x"46",x"DB",x"B4",x"D9",x"12",x"C2",x"3C", -- 0x0208
		x"FB",x"26",x"07",x"7A",x"6E",x"4B",x"10",x"09", -- 0x0210
		x"07",x"83",x"D2",x"FE",x"D2",x"7C",x"57",x"A1", -- 0x0218
		x"B1",x"4B",x"3C",x"75",x"AA",x"4A",x"9F",x"30", -- 0x0220
		x"90",x"7B",x"E5",x"6B",x"0D",x"A8",x"A7",x"88", -- 0x0228
		x"4E",x"2F",x"03",x"BC",x"F9",x"92",x"46",x"81", -- 0x0230
		x"95",x"19",x"80",x"68",x"15",x"58",x"0A",x"C6", -- 0x0238
		x"A3",x"C5",x"BC",x"CD",x"10",x"5C",x"FE",x"21", -- 0x0240
		x"57",x"64",x"8C",x"65",x"0D",x"B3",x"6D",x"DA", -- 0x0248
		x"E2",x"F0",x"98",x"5D",x"83",x"5E",x"DE",x"1A", -- 0x0250
		x"77",x"DE",x"82",x"8C",x"37",x"0D",x"D2",x"DB", -- 0x0258
		x"D2",x"8F",x"29",x"63",x"EB",x"28",x"84",x"C3", -- 0x0260
		x"8C",x"11",x"A8",x"19",x"C4",x"16",x"F4",x"28", -- 0x0268
		x"07",x"0D",x"85",x"0B",x"6B",x"E3",x"25",x"E2", -- 0x0270
		x"42",x"A7",x"EE",x"7A",x"B4",x"C1",x"D5",x"08", -- 0x0278
		x"D1",x"FE",x"6B",x"3D",x"A7",x"EF",x"01",x"34", -- 0x0280
		x"80",x"A9",x"CD",x"C4",x"40",x"C2",x"EC",x"47", -- 0x0288
		x"CF",x"F1",x"52",x"3B",x"55",x"F6",x"9D",x"98", -- 0x0290
		x"1F",x"0C",x"92",x"D3",x"CD",x"E7",x"5B",x"1F", -- 0x0298
		x"66",x"C6",x"5D",x"0E",x"36",x"DD",x"C2",x"B6", -- 0x02A0
		x"88",x"90",x"7C",x"C8",x"D2",x"E8",x"8F",x"A2", -- 0x02A8
		x"5B",x"62",x"5D",x"B0",x"59",x"7A",x"C8",x"78", -- 0x02B0
		x"86",x"5B",x"CC",x"D3",x"C2",x"28",x"F3",x"2A", -- 0x02B8
		x"6F",x"D0",x"38",x"A5",x"AE",x"7A",x"DC",x"B6", -- 0x02C0
		x"8A",x"59",x"FE",x"5D",x"C1",x"8F",x"7F",x"1D", -- 0x02C8
		x"F1",x"5C",x"4E",x"CA",x"D6",x"17",x"C3",x"5D", -- 0x02D0
		x"F2",x"90",x"32",x"35",x"38",x"26",x"5F",x"27", -- 0x02D8
		x"F6",x"18",x"CD",x"25",x"92",x"AA",x"DC",x"9D", -- 0x02E0
		x"83",x"DB",x"FA",x"45",x"EA",x"FA",x"E2",x"5C", -- 0x02E8
		x"57",x"B0",x"28",x"2F",x"C7",x"EB",x"8C",x"3A", -- 0x02F0
		x"FB",x"3E",x"70",x"34",x"64",x"4F",x"DB",x"DA", -- 0x02F8
		x"67",x"A9",x"01",x"7A",x"D3",x"5D",x"97",x"D6", -- 0x0300
		x"B8",x"92",x"9B",x"A4",x"0D",x"FD",x"01",x"65", -- 0x0308
		x"AE",x"A8",x"14",x"F6",x"14",x"20",x"31",x"10", -- 0x0310
		x"5F",x"21",x"C4",x"43",x"F0",x"A0",x"1F",x"58", -- 0x0318
		x"C9",x"9F",x"52",x"1D",x"7C",x"E9",x"F3",x"35", -- 0x0320
		x"FC",x"0F",x"D9",x"89",x"0E",x"5B",x"EE",x"BC", -- 0x0328
		x"04",x"82",x"B3",x"19",x"A3",x"65",x"A8",x"03", -- 0x0330
		x"06",x"6D",x"46",x"F6",x"8D",x"E4",x"CF",x"57", -- 0x0338
		x"04",x"22",x"74",x"80",x"8C",x"E7",x"B6",x"09", -- 0x0340
		x"77",x"10",x"92",x"85",x"EA",x"02",x"C1",x"EF", -- 0x0348
		x"84",x"76",x"88",x"28",x"5B",x"31",x"AA",x"61", -- 0x0350
		x"9F",x"71",x"59",x"AC",x"56",x"A8",x"05",x"DA", -- 0x0358
		x"4A",x"F8",x"5B",x"D6",x"61",x"91",x"5F",x"D8", -- 0x0360
		x"22",x"F2",x"DD",x"0D",x"74",x"9F",x"7C",x"F8", -- 0x0368
		x"95",x"05",x"A1",x"70",x"37",x"CB",x"D2",x"56", -- 0x0370
		x"BC",x"AB",x"03",x"93",x"54",x"87",x"6E",x"9E", -- 0x0378
		x"01",x"49",x"F5",x"62",x"DB",x"55",x"BA",x"7D", -- 0x0380
		x"C7",x"18",x"0A",x"BB",x"37",x"87",x"35",x"CD", -- 0x0388
		x"8C",x"56",x"BD",x"43",x"22",x"90",x"99",x"DF", -- 0x0390
		x"BB",x"1D",x"73",x"10",x"24",x"61",x"2F",x"25", -- 0x0398
		x"AA",x"25",x"87",x"06",x"F9",x"C1",x"83",x"42", -- 0x03A0
		x"D9",x"8E",x"FD",x"12",x"16",x"33",x"5F",x"22", -- 0x03A8
		x"09",x"1D",x"66",x"2C",x"2E",x"7F",x"8B",x"E9", -- 0x03B0
		x"1C",x"7E",x"7A",x"41",x"DF",x"29",x"66",x"8A", -- 0x03B8
		x"CD",x"6E",x"91",x"47",x"30",x"15",x"89",x"8A", -- 0x03C0
		x"23",x"08",x"1C",x"39",x"BA",x"7B",x"DB",x"C4", -- 0x03C8
		x"18",x"42",x"70",x"C5",x"41",x"FB",x"B0",x"5E", -- 0x03D0
		x"F9",x"AA",x"1F",x"D9",x"D3",x"85",x"E3",x"21", -- 0x03D8
		x"F3",x"75",x"68",x"A4",x"0B",x"72",x"AE",x"AD", -- 0x03E0
		x"7A",x"CA",x"67",x"B4",x"C5",x"43",x"F8",x"DD", -- 0x03E8
		x"05",x"69",x"A4",x"46",x"E4",x"D4",x"24",x"DE", -- 0x03F0
		x"FE",x"43",x"38",x"52",x"49",x"1D",x"73",x"BC", -- 0x03F8
		x"12",x"5B",x"61",x"9C",x"CD",x"8F",x"4B",x"C7", -- 0x0400
		x"5A",x"B2",x"7D",x"20",x"F5",x"76",x"7E",x"FA", -- 0x0408
		x"60",x"A2",x"C0",x"45",x"F6",x"E5",x"A4",x"75", -- 0x0410
		x"A8",x"5C",x"C7",x"F1",x"79",x"BA",x"AF",x"0C", -- 0x0418
		x"16",x"90",x"A8",x"64",x"21",x"73",x"2C",x"FA", -- 0x0420
		x"26",x"29",x"9B",x"9B",x"A0",x"99",x"96",x"01", -- 0x0428
		x"3C",x"D7",x"C5",x"B2",x"3D",x"E9",x"28",x"E5", -- 0x0430
		x"47",x"6F",x"58",x"40",x"A9",x"87",x"CB",x"3F", -- 0x0438
		x"97",x"75",x"A3",x"38",x"E8",x"D0",x"34",x"8F", -- 0x0440
		x"F9",x"4F",x"2B",x"1A",x"E8",x"42",x"9A",x"A4", -- 0x0448
		x"1A",x"E0",x"57",x"57",x"CA",x"FE",x"BC",x"91", -- 0x0450
		x"ED",x"94",x"D2",x"97",x"1C",x"9E",x"D6",x"B4", -- 0x0458
		x"93",x"7B",x"EC",x"FC",x"CB",x"A0",x"8C",x"45", -- 0x0460
		x"EF",x"37",x"DF",x"58",x"79",x"7A",x"FC",x"93", -- 0x0468
		x"5B",x"D3",x"6A",x"A6",x"52",x"28",x"38",x"40", -- 0x0470
		x"3C",x"0B",x"D7",x"59",x"2A",x"AF",x"8D",x"3D", -- 0x0478
		x"AA",x"F9",x"3A",x"F5",x"9B",x"46",x"3B",x"0B", -- 0x0480
		x"7E",x"9A",x"E3",x"F7",x"16",x"60",x"0C",x"F0", -- 0x0488
		x"35",x"76",x"17",x"07",x"1E",x"50",x"48",x"5B", -- 0x0490
		x"DA",x"9F",x"34",x"84",x"CE",x"C1",x"C2",x"79", -- 0x0498
		x"3B",x"FC",x"EE",x"D6",x"C3",x"AA",x"62",x"42", -- 0x04A0
		x"45",x"46",x"B9",x"DA",x"26",x"C5",x"CC",x"5B", -- 0x04A8
		x"BC",x"E3",x"E2",x"5A",x"B3",x"2B",x"B5",x"8F", -- 0x04B0
		x"4A",x"69",x"14",x"1A",x"AA",x"D6",x"13",x"E6", -- 0x04B8
		x"54",x"03",x"3D",x"18",x"AD",x"9F",x"D9",x"F2", -- 0x04C0
		x"65",x"93",x"4E",x"8C",x"D9",x"9A",x"67",x"16", -- 0x04C8
		x"7E",x"4A",x"70",x"B2",x"F4",x"A6",x"42",x"BF", -- 0x04D0
		x"10",x"D5",x"D9",x"BB",x"2D",x"EC",x"22",x"01", -- 0x04D8
		x"6F",x"5F",x"98",x"1D",x"7F",x"72",x"90",x"E4", -- 0x04E0
		x"85",x"5E",x"F0",x"DE",x"F8",x"D8",x"F4",x"77", -- 0x04E8
		x"23",x"66",x"A9",x"98",x"0D",x"6B",x"58",x"9C", -- 0x04F0
		x"42",x"B1",x"D7",x"EE",x"1E",x"F9",x"EF",x"8E", -- 0x04F8
		x"D9",x"88",x"2B",x"59",x"7A",x"3B",x"BD",x"7F", -- 0x0500
		x"99",x"AF",x"5F",x"92",x"88",x"54",x"8A",x"2B", -- 0x0508
		x"3A",x"34",x"43",x"C6",x"A0",x"1B",x"E3",x"62", -- 0x0510
		x"CC",x"BB",x"D0",x"6B",x"36",x"C0",x"F9",x"10", -- 0x0518
		x"C8",x"A4",x"69",x"43",x"E0",x"27",x"C2",x"F9", -- 0x0520
		x"56",x"A1",x"8D",x"5E",x"76",x"97",x"0A",x"B0", -- 0x0528
		x"4B",x"4D",x"F7",x"6B",x"69",x"DB",x"CD",x"B5", -- 0x0530
		x"17",x"9E",x"A0",x"4D",x"DE",x"9A",x"5D",x"A7", -- 0x0538
		x"BF",x"46",x"6A",x"A0",x"ED",x"AD",x"1A",x"C3", -- 0x0540
		x"4F",x"A7",x"23",x"C5",x"BE",x"2D",x"F6",x"0B", -- 0x0548
		x"7A",x"6E",x"76",x"63",x"4A",x"45",x"99",x"61", -- 0x0550
		x"63",x"3A",x"2F",x"C2",x"55",x"8C",x"E9",x"15", -- 0x0558
		x"53",x"D4",x"35",x"41",x"82",x"4F",x"05",x"51", -- 0x0560
		x"77",x"A7",x"97",x"36",x"D4",x"8E",x"41",x"CF", -- 0x0568
		x"7C",x"B8",x"B2",x"C6",x"7D",x"4C",x"A7",x"60", -- 0x0570
		x"07",x"D6",x"A2",x"DB",x"E3",x"8D",x"F0",x"37", -- 0x0578
		x"62",x"A5",x"F7",x"64",x"F4",x"7C",x"B5",x"EB", -- 0x0580
		x"25",x"4D",x"23",x"F9",x"5B",x"E3",x"49",x"D7", -- 0x0588
		x"9C",x"FC",x"1E",x"99",x"C8",x"46",x"7A",x"CF", -- 0x0590
		x"1D",x"1D",x"AB",x"80",x"AA",x"1C",x"37",x"8C", -- 0x0598
		x"C1",x"2F",x"F0",x"37",x"AC",x"A7",x"23",x"51", -- 0x05A0
		x"74",x"C5",x"CA",x"D0",x"AA",x"15",x"A8",x"C6", -- 0x05A8
		x"12",x"47",x"61",x"DA",x"8D",x"DB",x"2B",x"2A", -- 0x05B0
		x"78",x"56",x"AB",x"A3",x"73",x"E2",x"30",x"B4", -- 0x05B8
		x"92",x"A1",x"EB",x"BE",x"49",x"8F",x"10",x"BD", -- 0x05C0
		x"55",x"5A",x"0E",x"00",x"6F",x"37",x"C7",x"01", -- 0x05C8
		x"7E",x"A8",x"5C",x"0C",x"04",x"87",x"B5",x"7C", -- 0x05D0
		x"DD",x"E0",x"20",x"D0",x"C4",x"51",x"86",x"D6", -- 0x05D8
		x"72",x"F1",x"95",x"BB",x"81",x"25",x"F8",x"D7", -- 0x05E0
		x"7F",x"08",x"57",x"6F",x"3F",x"1F",x"70",x"3D", -- 0x05E8
		x"C7",x"CC",x"C8",x"CB",x"54",x"7E",x"C8",x"B2", -- 0x05F0
		x"60",x"E8",x"83",x"A4",x"B9",x"89",x"FA",x"2C", -- 0x05F8
		x"7C",x"10",x"67",x"FD",x"35",x"61",x"55",x"34", -- 0x0600
		x"E8",x"AD",x"A3",x"A7",x"4C",x"94",x"64",x"15", -- 0x0608
		x"61",x"2D",x"60",x"36",x"2B",x"29",x"68",x"0B", -- 0x0610
		x"92",x"EB",x"AF",x"4C",x"F5",x"AA",x"79",x"72", -- 0x0618
		x"BA",x"60",x"EF",x"6F",x"41",x"46",x"24",x"2A", -- 0x0620
		x"73",x"C7",x"51",x"BF",x"DB",x"B5",x"54",x"3E", -- 0x0628
		x"62",x"35",x"F3",x"8E",x"DD",x"5C",x"99",x"70", -- 0x0630
		x"C7",x"C9",x"BD",x"BD",x"F3",x"B6",x"AF",x"2F", -- 0x0638
		x"17",x"A0",x"9E",x"D8",x"66",x"42",x"82",x"59", -- 0x0640
		x"0B",x"D4",x"19",x"E6",x"0A",x"ED",x"A4",x"6D", -- 0x0648
		x"A2",x"98",x"7B",x"80",x"74",x"15",x"F1",x"3D", -- 0x0650
		x"5E",x"2F",x"7A",x"53",x"65",x"2B",x"82",x"FB", -- 0x0658
		x"4B",x"A0",x"D4",x"B1",x"E3",x"58",x"8A",x"6E", -- 0x0660
		x"AC",x"23",x"D4",x"B6",x"11",x"F9",x"A3",x"B3", -- 0x0668
		x"12",x"1F",x"B4",x"87",x"B4",x"26",x"44",x"13", -- 0x0670
		x"D4",x"BE",x"E5",x"3A",x"69",x"E7",x"B5",x"B4", -- 0x0678
		x"09",x"8B",x"E5",x"6C",x"63",x"70",x"5A",x"10", -- 0x0680
		x"94",x"2F",x"46",x"25",x"A8",x"EA",x"59",x"BB", -- 0x0688
		x"89",x"0E",x"C2",x"3E",x"34",x"07",x"D1",x"88", -- 0x0690
		x"45",x"B7",x"C2",x"AF",x"20",x"78",x"64",x"29", -- 0x0698
		x"83",x"CA",x"95",x"66",x"3B",x"EF",x"76",x"CF", -- 0x06A0
		x"9E",x"3D",x"F5",x"C7",x"A7",x"CE",x"83",x"31", -- 0x06A8
		x"DC",x"C5",x"EF",x"90",x"4C",x"41",x"19",x"91", -- 0x06B0
		x"78",x"5B",x"C0",x"98",x"53",x"A5",x"C1",x"D7", -- 0x06B8
		x"70",x"57",x"3E",x"AB",x"C6",x"35",x"FB",x"E5", -- 0x06C0
		x"F1",x"71",x"AD",x"99",x"40",x"31",x"4A",x"1D", -- 0x06C8
		x"76",x"B9",x"2D",x"C2",x"FA",x"46",x"D3",x"74", -- 0x06D0
		x"21",x"15",x"0D",x"74",x"BA",x"CF",x"4C",x"2B", -- 0x06D8
		x"A6",x"0B",x"56",x"ED",x"BF",x"52",x"D3",x"B1", -- 0x06E0
		x"43",x"81",x"CA",x"83",x"32",x"15",x"A0",x"A8", -- 0x06E8
		x"CF",x"4D",x"EA",x"4A",x"13",x"3E",x"BE",x"34", -- 0x06F0
		x"53",x"CC",x"A9",x"8D",x"1C",x"75",x"38",x"42", -- 0x06F8
		x"00",x"8F",x"30",x"BF",x"61",x"83",x"F0",x"A5", -- 0x0700
		x"05",x"BB",x"29",x"37",x"51",x"4A",x"5F",x"A0", -- 0x0708
		x"97",x"C9",x"EA",x"2B",x"09",x"2A",x"5F",x"DB", -- 0x0710
		x"76",x"88",x"6A",x"12",x"FE",x"A2",x"54",x"FE", -- 0x0718
		x"32",x"05",x"3F",x"14",x"88",x"30",x"B9",x"8E", -- 0x0720
		x"6C",x"62",x"45",x"3D",x"2C",x"25",x"DD",x"44", -- 0x0728
		x"EE",x"48",x"6F",x"F7",x"F1",x"CE",x"D4",x"68", -- 0x0730
		x"D7",x"BE",x"7A",x"D6",x"61",x"4F",x"55",x"14", -- 0x0738
		x"54",x"94",x"28",x"5C",x"C5",x"61",x"6A",x"B1", -- 0x0740
		x"C3",x"B0",x"EE",x"F0",x"55",x"4C",x"35",x"44", -- 0x0748
		x"14",x"24",x"BC",x"07",x"F2",x"11",x"EE",x"CA", -- 0x0750
		x"CF",x"E9",x"21",x"B0",x"39",x"77",x"C4",x"0D", -- 0x0758
		x"0C",x"EC",x"E8",x"51",x"CD",x"54",x"03",x"92", -- 0x0760
		x"84",x"71",x"03",x"D9",x"BD",x"B7",x"1E",x"D2", -- 0x0768
		x"DB",x"5A",x"59",x"4E",x"6B",x"C7",x"99",x"BA", -- 0x0770
		x"B1",x"BA",x"6C",x"6A",x"B1",x"31",x"F6",x"3E", -- 0x0778
		x"9E",x"E0",x"8F",x"6C",x"35",x"13",x"7E",x"B9", -- 0x0780
		x"84",x"81",x"13",x"C2",x"B8",x"31",x"15",x"94", -- 0x0788
		x"8C",x"6E",x"63",x"77",x"B5",x"FC",x"33",x"68", -- 0x0790
		x"37",x"9F",x"D2",x"E9",x"D0",x"4A",x"28",x"EE", -- 0x0798
		x"2B",x"37",x"5C",x"DF",x"C9",x"DA",x"99",x"CE", -- 0x07A0
		x"DC",x"AC",x"91",x"15",x"5D",x"A6",x"AA",x"69", -- 0x07A8
		x"94",x"0E",x"E1",x"4A",x"8A",x"94",x"32",x"C1", -- 0x07B0
		x"34",x"85",x"2B",x"84",x"CF",x"D2",x"74",x"7A", -- 0x07B8
		x"0B",x"50",x"5A",x"D4",x"2B",x"73",x"A3",x"87", -- 0x07C0
		x"20",x"B4",x"9D",x"FC",x"DA",x"C7",x"E6",x"EE", -- 0x07C8
		x"55",x"C8",x"B9",x"DF",x"5D",x"EB",x"21",x"11", -- 0x07D0
		x"71",x"4D",x"95",x"C0",x"9F",x"89",x"3B",x"AA", -- 0x07D8
		x"D9",x"95",x"00",x"85",x"09",x"23",x"0D",x"A8", -- 0x07E0
		x"58",x"2A",x"26",x"33",x"F1",x"0D",x"23",x"C6", -- 0x07E8
		x"55",x"DC",x"26",x"32",x"48",x"48",x"43",x"3A", -- 0x07F0
		x"15",x"58",x"7A",x"B4",x"62",x"B6",x"DF",x"3C", -- 0x07F8
		x"CB",x"5F",x"41",x"55",x"82",x"4F",x"7D",x"DA", -- 0x0800
		x"F8",x"A3",x"8E",x"6B",x"30",x"31",x"32",x"85", -- 0x0808
		x"8D",x"59",x"B7",x"D5",x"21",x"7A",x"8F",x"B5", -- 0x0810
		x"53",x"0B",x"6A",x"B5",x"41",x"C9",x"71",x"0D", -- 0x0818
		x"29",x"B3",x"62",x"2C",x"82",x"60",x"07",x"7B", -- 0x0820
		x"04",x"15",x"66",x"35",x"46",x"19",x"3A",x"D3", -- 0x0828
		x"72",x"F2",x"2A",x"13",x"EC",x"39",x"C8",x"40", -- 0x0830
		x"44",x"B2",x"75",x"85",x"7D",x"67",x"13",x"26", -- 0x0838
		x"1B",x"75",x"52",x"9D",x"D5",x"D9",x"98",x"5A", -- 0x0840
		x"EE",x"7F",x"0F",x"B5",x"98",x"49",x"09",x"8A", -- 0x0848
		x"BB",x"33",x"9D",x"A9",x"EC",x"E5",x"69",x"31", -- 0x0850
		x"98",x"5F",x"37",x"95",x"C6",x"4A",x"BC",x"E1", -- 0x0858
		x"3F",x"0F",x"FE",x"95",x"E8",x"17",x"EF",x"58", -- 0x0860
		x"96",x"7E",x"0E",x"2F",x"C7",x"17",x"B9",x"84", -- 0x0868
		x"CA",x"D6",x"AD",x"B7",x"BC",x"96",x"68",x"D5", -- 0x0870
		x"F5",x"9F",x"6B",x"3C",x"E9",x"A7",x"9D",x"2A", -- 0x0878
		x"B7",x"9C",x"BF",x"20",x"34",x"2F",x"78",x"CA", -- 0x0880
		x"AD",x"86",x"FA",x"F4",x"9E",x"34",x"79",x"E8", -- 0x0888
		x"0C",x"A6",x"A0",x"48",x"3E",x"88",x"1E",x"B3", -- 0x0890
		x"29",x"8A",x"F0",x"13",x"32",x"8E",x"BC",x"69", -- 0x0898
		x"AB",x"FB",x"8A",x"DF",x"AA",x"03",x"AA",x"58", -- 0x08A0
		x"0A",x"25",x"4E",x"28",x"D9",x"47",x"11",x"E5", -- 0x08A8
		x"6E",x"31",x"2E",x"AC",x"B9",x"CC",x"DF",x"E2", -- 0x08B0
		x"57",x"D0",x"76",x"09",x"DF",x"B2",x"F2",x"8B", -- 0x08B8
		x"AF",x"FC",x"EA",x"D9",x"7F",x"15",x"33",x"89", -- 0x08C0
		x"3B",x"01",x"B1",x"15",x"C7",x"42",x"7A",x"36", -- 0x08C8
		x"73",x"28",x"62",x"AD",x"F4",x"43",x"10",x"CB", -- 0x08D0
		x"93",x"06",x"55",x"73",x"B9",x"48",x"7E",x"E8", -- 0x08D8
		x"45",x"69",x"C2",x"C4",x"7F",x"75",x"CE",x"3A", -- 0x08E0
		x"F5",x"00",x"CE",x"BE",x"43",x"C8",x"74",x"36", -- 0x08E8
		x"F0",x"57",x"E3",x"66",x"9A",x"F4",x"32",x"2E", -- 0x08F0
		x"FA",x"07",x"22",x"B4",x"4F",x"A0",x"1D",x"14", -- 0x08F8
		x"0B",x"E0",x"59",x"0A",x"D5",x"28",x"C3",x"CC", -- 0x0900
		x"28",x"12",x"0B",x"EA",x"DA",x"FE",x"22",x"4B", -- 0x0908
		x"56",x"06",x"B1",x"F0",x"7A",x"64",x"9F",x"76", -- 0x0910
		x"6B",x"C1",x"AA",x"3B",x"62",x"C8",x"4F",x"EC", -- 0x0918
		x"29",x"28",x"76",x"FE",x"CF",x"3A",x"4B",x"78", -- 0x0920
		x"4C",x"56",x"63",x"27",x"56",x"85",x"F2",x"AC", -- 0x0928
		x"0C",x"A4",x"1E",x"86",x"09",x"BD",x"FC",x"F4", -- 0x0930
		x"7F",x"28",x"30",x"E1",x"70",x"7F",x"4F",x"99", -- 0x0938
		x"28",x"C5",x"18",x"F7",x"80",x"E3",x"70",x"CC", -- 0x0940
		x"3A",x"54",x"74",x"10",x"D9",x"67",x"3D",x"E5", -- 0x0948
		x"8B",x"5B",x"EC",x"15",x"19",x"E9",x"0A",x"18", -- 0x0950
		x"91",x"3A",x"79",x"02",x"39",x"C8",x"1B",x"61", -- 0x0958
		x"0F",x"B3",x"5A",x"8F",x"97",x"4A",x"DB",x"D1", -- 0x0960
		x"9E",x"50",x"62",x"F8",x"37",x"9F",x"5E",x"43", -- 0x0968
		x"7A",x"4B",x"58",x"13",x"B5",x"E1",x"2B",x"47", -- 0x0970
		x"1C",x"A4",x"C9",x"D4",x"ED",x"E4",x"37",x"FC", -- 0x0978
		x"98",x"11",x"8C",x"AF",x"DA",x"68",x"02",x"7A", -- 0x0980
		x"39",x"64",x"F2",x"EF",x"83",x"51",x"33",x"FD", -- 0x0988
		x"1D",x"0B",x"11",x"D2",x"EC",x"3C",x"99",x"88", -- 0x0990
		x"60",x"63",x"5E",x"4E",x"C8",x"95",x"4B",x"E0", -- 0x0998
		x"26",x"57",x"91",x"01",x"C0",x"93",x"FA",x"79", -- 0x09A0
		x"77",x"6D",x"69",x"FA",x"3F",x"1D",x"78",x"5C", -- 0x09A8
		x"A7",x"89",x"AE",x"95",x"45",x"48",x"1E",x"25", -- 0x09B0
		x"2C",x"FB",x"74",x"F4",x"91",x"3F",x"D5",x"37", -- 0x09B8
		x"97",x"E6",x"B8",x"D7",x"F9",x"B3",x"51",x"71", -- 0x09C0
		x"A1",x"3A",x"EB",x"E0",x"D6",x"64",x"3D",x"7F", -- 0x09C8
		x"6D",x"EB",x"15",x"32",x"34",x"B2",x"58",x"DF", -- 0x09D0
		x"AF",x"4C",x"D4",x"C0",x"8B",x"2B",x"78",x"23", -- 0x09D8
		x"12",x"31",x"7A",x"0D",x"64",x"4B",x"7E",x"06", -- 0x09E0
		x"86",x"EA",x"E6",x"5D",x"4F",x"24",x"5C",x"3D", -- 0x09E8
		x"8F",x"71",x"6F",x"44",x"A4",x"C7",x"24",x"D3", -- 0x09F0
		x"14",x"F9",x"14",x"20",x"A4",x"8C",x"C2",x"B6", -- 0x09F8
		x"BD",x"3E",x"C3",x"23",x"89",x"C2",x"A8",x"8F", -- 0x0A00
		x"AD",x"90",x"6D",x"7C",x"34",x"C9",x"B9",x"44", -- 0x0A08
		x"BB",x"A9",x"88",x"DF",x"71",x"AC",x"B3",x"06", -- 0x0A10
		x"26",x"C7",x"A5",x"CA",x"D4",x"68",x"02",x"92", -- 0x0A18
		x"26",x"45",x"35",x"30",x"87",x"DE",x"3F",x"35", -- 0x0A20
		x"EE",x"AC",x"32",x"A2",x"F6",x"6B",x"E6",x"B2", -- 0x0A28
		x"15",x"6F",x"12",x"07",x"9C",x"C5",x"8C",x"42", -- 0x0A30
		x"0D",x"32",x"8D",x"E1",x"1A",x"8F",x"F4",x"41", -- 0x0A38
		x"D4",x"A9",x"F0",x"5D",x"08",x"30",x"12",x"F6", -- 0x0A40
		x"DD",x"C3",x"1A",x"54",x"30",x"01",x"07",x"45", -- 0x0A48
		x"F0",x"98",x"CB",x"0D",x"DD",x"58",x"4F",x"EA", -- 0x0A50
		x"0A",x"DC",x"4D",x"25",x"6C",x"C1",x"E5",x"C1", -- 0x0A58
		x"6B",x"D6",x"1F",x"74",x"86",x"B0",x"EA",x"64", -- 0x0A60
		x"75",x"05",x"B8",x"A5",x"86",x"3F",x"6A",x"77", -- 0x0A68
		x"57",x"37",x"84",x"35",x"0F",x"53",x"A0",x"1A", -- 0x0A70
		x"31",x"6D",x"BE",x"1D",x"2F",x"A4",x"DE",x"9A", -- 0x0A78
		x"FA",x"FD",x"8E",x"81",x"AF",x"7A",x"66",x"A4", -- 0x0A80
		x"7F",x"9E",x"4A",x"85",x"5E",x"34",x"FC",x"B5", -- 0x0A88
		x"EA",x"01",x"6B",x"FA",x"55",x"0C",x"94",x"06", -- 0x0A90
		x"79",x"53",x"23",x"A8",x"77",x"82",x"C2",x"F1", -- 0x0A98
		x"00",x"52",x"73",x"2F",x"CC",x"59",x"D3",x"CB", -- 0x0AA0
		x"F8",x"1E",x"52",x"D6",x"D2",x"CE",x"0C",x"BD", -- 0x0AA8
		x"50",x"77",x"B8",x"25",x"83",x"4D",x"AA",x"7C", -- 0x0AB0
		x"20",x"CD",x"25",x"97",x"CF",x"E8",x"89",x"D0", -- 0x0AB8
		x"BA",x"7D",x"00",x"87",x"D6",x"54",x"D2",x"4F", -- 0x0AC0
		x"F1",x"A4",x"26",x"C4",x"74",x"33",x"83",x"44", -- 0x0AC8
		x"2A",x"3C",x"69",x"AE",x"0A",x"14",x"2B",x"A9", -- 0x0AD0
		x"61",x"D0",x"C1",x"32",x"39",x"CA",x"82",x"F3", -- 0x0AD8
		x"48",x"02",x"FA",x"9F",x"56",x"CD",x"6E",x"49", -- 0x0AE0
		x"73",x"95",x"0E",x"67",x"48",x"91",x"AB",x"72", -- 0x0AE8
		x"4E",x"15",x"A0",x"D7",x"A8",x"CC",x"81",x"0A", -- 0x0AF0
		x"1D",x"43",x"BB",x"56",x"0F",x"3E",x"4A",x"D6", -- 0x0AF8
		x"41",x"45",x"76",x"17",x"92",x"E5",x"60",x"85", -- 0x0B00
		x"FA",x"EE",x"EC",x"C2",x"80",x"98",x"B4",x"4E", -- 0x0B08
		x"2D",x"56",x"26",x"55",x"A2",x"A8",x"60",x"BF", -- 0x0B10
		x"EB",x"9B",x"95",x"7A",x"5A",x"5F",x"52",x"1B", -- 0x0B18
		x"24",x"48",x"32",x"B6",x"AD",x"93",x"3D",x"28", -- 0x0B20
		x"82",x"A9",x"6A",x"82",x"43",x"20",x"D1",x"EF", -- 0x0B28
		x"F5",x"F7",x"46",x"18",x"20",x"26",x"D7",x"8C", -- 0x0B30
		x"C1",x"EC",x"07",x"1C",x"4C",x"D8",x"37",x"70", -- 0x0B38
		x"A1",x"E9",x"A6",x"CE",x"FC",x"E3",x"77",x"FE", -- 0x0B40
		x"8E",x"E1",x"81",x"51",x"81",x"D2",x"C0",x"77", -- 0x0B48
		x"4B",x"07",x"8F",x"6B",x"AC",x"E6",x"F7",x"6F", -- 0x0B50
		x"53",x"7F",x"0B",x"9F",x"D7",x"C2",x"8F",x"F8", -- 0x0B58
		x"2C",x"37",x"48",x"29",x"9A",x"BF",x"28",x"29", -- 0x0B60
		x"21",x"29",x"F9",x"A3",x"7C",x"BB",x"9A",x"C7", -- 0x0B68
		x"42",x"AA",x"B2",x"EF",x"11",x"2B",x"DE",x"65", -- 0x0B70
		x"2A",x"69",x"05",x"81",x"AB",x"15",x"7B",x"D7", -- 0x0B78
		x"4C",x"C3",x"80",x"E6",x"03",x"A8",x"90",x"24", -- 0x0B80
		x"52",x"8A",x"47",x"CE",x"C5",x"E2",x"16",x"88", -- 0x0B88
		x"0D",x"C8",x"F7",x"1E",x"73",x"56",x"83",x"9D", -- 0x0B90
		x"BF",x"09",x"20",x"EB",x"1E",x"1B",x"C3",x"E9", -- 0x0B98
		x"5E",x"45",x"D0",x"61",x"6D",x"61",x"85",x"3F", -- 0x0BA0
		x"6C",x"CD",x"0E",x"32",x"30",x"A3",x"3A",x"3D", -- 0x0BA8
		x"EC",x"32",x"DA",x"60",x"88",x"DE",x"7E",x"C8", -- 0x0BB0
		x"67",x"9E",x"B4",x"85",x"B9",x"F7",x"6F",x"18", -- 0x0BB8
		x"BC",x"BF",x"F8",x"2B",x"22",x"7E",x"E9",x"0E", -- 0x0BC0
		x"CB",x"F8",x"BF",x"7B",x"1C",x"FA",x"38",x"09", -- 0x0BC8
		x"2D",x"93",x"6A",x"36",x"72",x"E8",x"FE",x"D9", -- 0x0BD0
		x"07",x"33",x"DE",x"40",x"2B",x"CD",x"D7",x"68", -- 0x0BD8
		x"8D",x"D0",x"13",x"2F",x"CE",x"FC",x"3D",x"1B", -- 0x0BE0
		x"F5",x"FD",x"16",x"92",x"F8",x"4F",x"9B",x"A5", -- 0x0BE8
		x"E2",x"06",x"DB",x"D4",x"6E",x"DA",x"AE",x"75", -- 0x0BF0
		x"8D",x"8D",x"35",x"B9",x"5B",x"0D",x"22",x"68", -- 0x0BF8
		x"DD",x"35",x"98",x"2D",x"32",x"D5",x"48",x"A8", -- 0x0C00
		x"53",x"5E",x"3B",x"CB",x"2D",x"56",x"72",x"8F", -- 0x0C08
		x"DC",x"4E",x"64",x"4B",x"A9",x"92",x"41",x"37", -- 0x0C10
		x"20",x"F5",x"70",x"FA",x"04",x"12",x"64",x"61", -- 0x0C18
		x"C6",x"7C",x"8E",x"F9",x"D1",x"56",x"22",x"26", -- 0x0C20
		x"35",x"DC",x"F1",x"62",x"33",x"64",x"72",x"10", -- 0x0C28
		x"33",x"D6",x"DB",x"5C",x"E9",x"9C",x"93",x"0A", -- 0x0C30
		x"92",x"84",x"85",x"96",x"96",x"69",x"78",x"5E", -- 0x0C38
		x"E5",x"07",x"D7",x"B7",x"DD",x"F9",x"5D",x"13", -- 0x0C40
		x"56",x"50",x"75",x"09",x"34",x"E7",x"99",x"E6", -- 0x0C48
		x"3F",x"75",x"43",x"29",x"91",x"D7",x"B2",x"24", -- 0x0C50
		x"5C",x"B7",x"3B",x"72",x"A0",x"B3",x"D0",x"86", -- 0x0C58
		x"3A",x"A8",x"BE",x"18",x"22",x"1C",x"2B",x"F7", -- 0x0C60
		x"EB",x"21",x"02",x"A0",x"88",x"9B",x"87",x"47", -- 0x0C68
		x"90",x"CB",x"EF",x"22",x"23",x"23",x"C5",x"FE", -- 0x0C70
		x"DA",x"01",x"F0",x"7C",x"34",x"C2",x"82",x"EE", -- 0x0C78
		x"EA",x"C0",x"07",x"8D",x"5D",x"B2",x"85",x"C8", -- 0x0C80
		x"53",x"07",x"69",x"DB",x"A2",x"71",x"A3",x"B2", -- 0x0C88
		x"BC",x"93",x"54",x"5F",x"B6",x"1B",x"DD",x"12", -- 0x0C90
		x"9B",x"CE",x"0E",x"50",x"91",x"10",x"3F",x"FC", -- 0x0C98
		x"D1",x"C5",x"8A",x"2F",x"78",x"8F",x"F7",x"4B", -- 0x0CA0
		x"97",x"E1",x"28",x"B9",x"53",x"CB",x"EC",x"8F", -- 0x0CA8
		x"DE",x"41",x"EE",x"96",x"DB",x"CC",x"28",x"78", -- 0x0CB0
		x"9B",x"36",x"48",x"AD",x"C5",x"87",x"AA",x"97", -- 0x0CB8
		x"4D",x"B4",x"46",x"46",x"44",x"BE",x"91",x"5B", -- 0x0CC0
		x"A0",x"39",x"16",x"73",x"84",x"03",x"82",x"64", -- 0x0CC8
		x"C3",x"71",x"FA",x"A0",x"BD",x"A2",x"98",x"59", -- 0x0CD0
		x"58",x"E0",x"86",x"1E",x"68",x"B0",x"36",x"35", -- 0x0CD8
		x"65",x"7C",x"FA",x"2A",x"BA",x"0D",x"85",x"DA", -- 0x0CE0
		x"46",x"1B",x"4E",x"CB",x"9D",x"50",x"AF",x"62", -- 0x0CE8
		x"C1",x"2A",x"82",x"7F",x"CC",x"1B",x"59",x"25", -- 0x0CF0
		x"FB",x"DF",x"C2",x"E3",x"11",x"F8",x"98",x"76", -- 0x0CF8
		x"F5",x"94",x"A0",x"30",x"21",x"A6",x"0C",x"E6", -- 0x0D00
		x"41",x"D9",x"32",x"DF",x"2B",x"E1",x"C1",x"EC", -- 0x0D08
		x"0C",x"44",x"EC",x"D8",x"DE",x"C5",x"7D",x"5A", -- 0x0D10
		x"25",x"C0",x"3E",x"36",x"39",x"56",x"2D",x"AE", -- 0x0D18
		x"EA",x"4D",x"DF",x"8B",x"F3",x"EB",x"73",x"36", -- 0x0D20
		x"C5",x"A5",x"95",x"F0",x"88",x"D6",x"5E",x"14", -- 0x0D28
		x"1B",x"CA",x"ED",x"79",x"90",x"EA",x"D3",x"35", -- 0x0D30
		x"AB",x"12",x"6C",x"65",x"68",x"99",x"14",x"D3", -- 0x0D38
		x"66",x"F3",x"DE",x"5B",x"DF",x"52",x"11",x"26", -- 0x0D40
		x"F8",x"26",x"96",x"01",x"FC",x"74",x"15",x"97", -- 0x0D48
		x"3F",x"82",x"11",x"4F",x"ED",x"E4",x"85",x"19", -- 0x0D50
		x"76",x"71",x"7E",x"5E",x"8A",x"93",x"B1",x"F0", -- 0x0D58
		x"07",x"91",x"CB",x"67",x"E3",x"5C",x"8D",x"5C", -- 0x0D60
		x"82",x"24",x"DC",x"7F",x"19",x"F2",x"96",x"58", -- 0x0D68
		x"F4",x"A7",x"28",x"E2",x"0C",x"AD",x"FC",x"02", -- 0x0D70
		x"9E",x"FA",x"61",x"A8",x"8E",x"92",x"19",x"16", -- 0x0D78
		x"24",x"E5",x"7D",x"88",x"42",x"0B",x"E4",x"C5", -- 0x0D80
		x"AE",x"42",x"C4",x"C7",x"B4",x"5C",x"A0",x"A9", -- 0x0D88
		x"83",x"C8",x"0D",x"10",x"F5",x"0A",x"12",x"14", -- 0x0D90
		x"05",x"F2",x"BC",x"14",x"86",x"D5",x"2A",x"AA", -- 0x0D98
		x"BB",x"27",x"33",x"7E",x"B1",x"98",x"C3",x"60", -- 0x0DA0
		x"DA",x"08",x"A8",x"0F",x"E3",x"C8",x"B8",x"68", -- 0x0DA8
		x"91",x"C5",x"F7",x"07",x"4F",x"0A",x"1B",x"D4", -- 0x0DB0
		x"FD",x"D7",x"E8",x"84",x"AD",x"92",x"AE",x"E9", -- 0x0DB8
		x"B9",x"62",x"E7",x"6B",x"FA",x"AB",x"4B",x"55", -- 0x0DC0
		x"B3",x"73",x"64",x"18",x"3C",x"9C",x"80",x"4D", -- 0x0DC8
		x"63",x"78",x"54",x"32",x"02",x"EE",x"07",x"00", -- 0x0DD0
		x"C6",x"6F",x"04",x"F4",x"81",x"B3",x"5E",x"3B", -- 0x0DD8
		x"95",x"46",x"26",x"90",x"71",x"F1",x"65",x"A4", -- 0x0DE0
		x"E4",x"49",x"BC",x"A1",x"65",x"BC",x"EE",x"48", -- 0x0DE8
		x"B4",x"C3",x"7B",x"B7",x"B2",x"82",x"37",x"F9", -- 0x0DF0
		x"72",x"BB",x"6E",x"F3",x"EE",x"CC",x"AF",x"84", -- 0x0DF8
		x"92",x"D5",x"94",x"83",x"47",x"79",x"28",x"2D", -- 0x0E00
		x"C2",x"65",x"CE",x"A7",x"A1",x"3D",x"F0",x"D6", -- 0x0E08
		x"80",x"6C",x"8E",x"B3",x"6E",x"45",x"2D",x"E0", -- 0x0E10
		x"80",x"9B",x"D5",x"6F",x"E7",x"85",x"F3",x"7A", -- 0x0E18
		x"DA",x"88",x"FD",x"23",x"02",x"A5",x"CF",x"44", -- 0x0E20
		x"8A",x"1E",x"EC",x"2D",x"5B",x"5D",x"04",x"5C", -- 0x0E28
		x"49",x"12",x"8F",x"B7",x"D6",x"BC",x"19",x"58", -- 0x0E30
		x"58",x"6E",x"47",x"40",x"F3",x"3C",x"3A",x"4E", -- 0x0E38
		x"44",x"B7",x"F0",x"C6",x"5D",x"C0",x"8A",x"68", -- 0x0E40
		x"DE",x"F6",x"15",x"BA",x"54",x"19",x"17",x"9D", -- 0x0E48
		x"AA",x"A6",x"56",x"01",x"E2",x"EE",x"59",x"3B", -- 0x0E50
		x"5D",x"21",x"FA",x"D0",x"5D",x"35",x"1F",x"21", -- 0x0E58
		x"6C",x"11",x"E7",x"C9",x"51",x"F2",x"B1",x"31", -- 0x0E60
		x"E9",x"C6",x"6B",x"3F",x"5F",x"02",x"5C",x"89", -- 0x0E68
		x"A8",x"32",x"8B",x"0B",x"21",x"64",x"46",x"7E", -- 0x0E70
		x"85",x"C0",x"4F",x"62",x"75",x"EE",x"84",x"E1", -- 0x0E78
		x"00",x"EB",x"2B",x"D0",x"DE",x"DD",x"81",x"49", -- 0x0E80
		x"A4",x"EC",x"88",x"84",x"EE",x"64",x"0E",x"17", -- 0x0E88
		x"97",x"99",x"22",x"B8",x"7E",x"E7",x"B7",x"04", -- 0x0E90
		x"A8",x"07",x"67",x"1E",x"75",x"6B",x"00",x"F4", -- 0x0E98
		x"D6",x"2C",x"C6",x"36",x"89",x"48",x"7F",x"2E", -- 0x0EA0
		x"36",x"87",x"32",x"A4",x"EB",x"41",x"BC",x"83", -- 0x0EA8
		x"5A",x"5E",x"BC",x"D8",x"47",x"74",x"DD",x"EF", -- 0x0EB0
		x"FA",x"C4",x"8E",x"71",x"AF",x"0E",x"E5",x"86", -- 0x0EB8
		x"3A",x"AC",x"BC",x"C3",x"F5",x"BB",x"72",x"AB", -- 0x0EC0
		x"43",x"A4",x"CF",x"AF",x"65",x"8C",x"33",x"C0", -- 0x0EC8
		x"6B",x"6F",x"19",x"B2",x"63",x"F6",x"22",x"5F", -- 0x0ED0
		x"3B",x"30",x"50",x"EA",x"3F",x"36",x"72",x"79", -- 0x0ED8
		x"63",x"AE",x"BD",x"D8",x"6B",x"AF",x"84",x"AE", -- 0x0EE0
		x"D3",x"54",x"5E",x"3A",x"61",x"12",x"7A",x"4C", -- 0x0EE8
		x"01",x"93",x"FE",x"65",x"0B",x"A0",x"44",x"46", -- 0x0EF0
		x"D1",x"94",x"B1",x"11",x"4A",x"24",x"0A",x"AD", -- 0x0EF8
		x"52",x"47",x"86",x"BD",x"F6",x"8A",x"EC",x"CB", -- 0x0F00
		x"5F",x"CA",x"85",x"40",x"DC",x"7F",x"8C",x"5E", -- 0x0F08
		x"92",x"0B",x"C3",x"9D",x"2B",x"08",x"64",x"FC", -- 0x0F10
		x"1C",x"16",x"8D",x"E5",x"B9",x"18",x"94",x"0C", -- 0x0F18
		x"5F",x"9A",x"CA",x"D6",x"A5",x"37",x"22",x"05", -- 0x0F20
		x"02",x"27",x"C4",x"5F",x"A6",x"D0",x"BD",x"39", -- 0x0F28
		x"5B",x"81",x"57",x"86",x"09",x"BB",x"04",x"25", -- 0x0F30
		x"51",x"11",x"0B",x"0B",x"29",x"1F",x"96",x"09", -- 0x0F38
		x"3A",x"E0",x"5F",x"DF",x"18",x"81",x"64",x"1B", -- 0x0F40
		x"28",x"A8",x"7A",x"4E",x"79",x"B7",x"87",x"D4", -- 0x0F48
		x"39",x"5E",x"5B",x"C1",x"99",x"DE",x"66",x"EA", -- 0x0F50
		x"F0",x"71",x"75",x"1A",x"11",x"8C",x"A2",x"CA", -- 0x0F58
		x"6D",x"02",x"AA",x"06",x"03",x"8E",x"A0",x"2B", -- 0x0F60
		x"37",x"9A",x"79",x"30",x"52",x"81",x"05",x"0B", -- 0x0F68
		x"5F",x"DF",x"CC",x"F9",x"BF",x"33",x"64",x"B0", -- 0x0F70
		x"24",x"5A",x"4A",x"B4",x"E6",x"ED",x"7F",x"D3", -- 0x0F78
		x"6F",x"2A",x"D9",x"73",x"38",x"7A",x"1E",x"6F", -- 0x0F80
		x"15",x"18",x"1F",x"67",x"19",x"24",x"F1",x"78", -- 0x0F88
		x"84",x"BE",x"F1",x"44",x"71",x"D6",x"74",x"96", -- 0x0F90
		x"31",x"3E",x"4B",x"97",x"2C",x"CB",x"6B",x"1C", -- 0x0F98
		x"75",x"46",x"0F",x"AE",x"40",x"2D",x"9D",x"D5", -- 0x0FA0
		x"C4",x"BD",x"BC",x"5D",x"61",x"AF",x"D6",x"E5", -- 0x0FA8
		x"6E",x"48",x"A9",x"60",x"1F",x"9D",x"F6",x"CF", -- 0x0FB0
		x"DC",x"C1",x"67",x"88",x"8D",x"53",x"A4",x"83", -- 0x0FB8
		x"99",x"B3",x"B1",x"59",x"61",x"4F",x"2F",x"26", -- 0x0FC0
		x"8C",x"EC",x"84",x"EE",x"1C",x"DA",x"54",x"0A", -- 0x0FC8
		x"A2",x"7E",x"6A",x"42",x"9B",x"61",x"12",x"78", -- 0x0FD0
		x"24",x"F9",x"02",x"31",x"4D",x"26",x"B4",x"66", -- 0x0FD8
		x"DA",x"66",x"BF",x"3C",x"36",x"EF",x"E1",x"C2", -- 0x0FE0
		x"5C",x"E5",x"31",x"78",x"C0",x"06",x"82",x"64", -- 0x0FE8
		x"04",x"ED",x"A6",x"9F",x"CE",x"38",x"19",x"72", -- 0x0FF0
		x"32",x"9A",x"A4",x"7F",x"C0",x"D8",x"E5",x"1B", -- 0x0FF8
		x"BF",x"A6",x"57",x"F5",x"16",x"B9",x"38",x"F1", -- 0x1000
		x"9F",x"E9",x"E9",x"61",x"EF",x"EB",x"45",x"F3", -- 0x1008
		x"59",x"6B",x"93",x"29",x"A3",x"2C",x"1B",x"56", -- 0x1010
		x"C6",x"3F",x"D5",x"08",x"19",x"3C",x"23",x"58", -- 0x1018
		x"E2",x"FA",x"CD",x"78",x"B4",x"06",x"E9",x"54", -- 0x1020
		x"EF",x"D3",x"35",x"5F",x"BF",x"F9",x"53",x"99", -- 0x1028
		x"E4",x"67",x"C2",x"89",x"93",x"5D",x"DF",x"DA", -- 0x1030
		x"9D",x"35",x"62",x"36",x"71",x"85",x"8E",x"D3", -- 0x1038
		x"00",x"5C",x"CB",x"B4",x"E1",x"B5",x"89",x"52", -- 0x1040
		x"09",x"3E",x"B1",x"49",x"B8",x"85",x"E2",x"9D", -- 0x1048
		x"6C",x"25",x"27",x"7F",x"82",x"86",x"D9",x"9F", -- 0x1050
		x"3C",x"3C",x"D5",x"2D",x"C2",x"E3",x"02",x"C2", -- 0x1058
		x"BF",x"4D",x"F7",x"A2",x"04",x"01",x"F4",x"8C", -- 0x1060
		x"BE",x"26",x"55",x"77",x"2B",x"38",x"16",x"97", -- 0x1068
		x"DC",x"BC",x"97",x"DF",x"C3",x"71",x"7F",x"00", -- 0x1070
		x"AE",x"D5",x"2D",x"F0",x"B9",x"AE",x"33",x"7A", -- 0x1078
		x"FC",x"2B",x"9C",x"80",x"AB",x"11",x"0D",x"6B", -- 0x1080
		x"37",x"63",x"E2",x"E2",x"1B",x"F8",x"F9",x"F8", -- 0x1088
		x"36",x"91",x"D8",x"F9",x"04",x"D7",x"79",x"B2", -- 0x1090
		x"AD",x"A6",x"A3",x"E7",x"D5",x"D6",x"E1",x"D2", -- 0x1098
		x"82",x"7E",x"53",x"AD",x"8F",x"DF",x"19",x"46", -- 0x10A0
		x"43",x"7C",x"A8",x"DE",x"F4",x"A3",x"D7",x"2B", -- 0x10A8
		x"35",x"30",x"25",x"39",x"87",x"1E",x"EB",x"B5", -- 0x10B0
		x"C5",x"0F",x"9D",x"9B",x"E6",x"7F",x"ED",x"E8", -- 0x10B8
		x"7D",x"41",x"96",x"8C",x"21",x"B0",x"D2",x"E4", -- 0x10C0
		x"AC",x"7C",x"C3",x"A1",x"9F",x"1B",x"CD",x"D4", -- 0x10C8
		x"CA",x"72",x"0F",x"52",x"91",x"7A",x"08",x"D6", -- 0x10D0
		x"8A",x"25",x"F1",x"F0",x"A4",x"DF",x"D9",x"22", -- 0x10D8
		x"A0",x"70",x"2E",x"41",x"A0",x"02",x"26",x"4D", -- 0x10E0
		x"FD",x"69",x"6F",x"1D",x"04",x"3D",x"F1",x"CE", -- 0x10E8
		x"2F",x"01",x"A1",x"C0",x"7C",x"A9",x"17",x"86", -- 0x10F0
		x"4F",x"09",x"77",x"F3",x"68",x"51",x"96",x"09", -- 0x10F8
		x"41",x"C4",x"CA",x"62",x"46",x"F0",x"AF",x"C3", -- 0x1100
		x"DA",x"1F",x"E0",x"DE",x"DB",x"D3",x"2E",x"0C", -- 0x1108
		x"54",x"CF",x"4C",x"50",x"F8",x"E3",x"D6",x"48", -- 0x1110
		x"EC",x"4E",x"BC",x"D5",x"9F",x"53",x"5E",x"61", -- 0x1118
		x"97",x"29",x"C3",x"5E",x"9A",x"F2",x"22",x"75", -- 0x1120
		x"13",x"83",x"D3",x"6E",x"D6",x"02",x"F9",x"2B", -- 0x1128
		x"D1",x"C6",x"7C",x"4B",x"AA",x"D2",x"93",x"17", -- 0x1130
		x"22",x"CF",x"EC",x"41",x"23",x"4C",x"A2",x"3B", -- 0x1138
		x"75",x"66",x"99",x"10",x"5A",x"3B",x"05",x"EC", -- 0x1140
		x"BE",x"D9",x"DA",x"15",x"5B",x"D5",x"41",x"AD", -- 0x1148
		x"9C",x"3D",x"F8",x"C6",x"10",x"0C",x"DD",x"B1", -- 0x1150
		x"DC",x"4B",x"F3",x"7F",x"97",x"16",x"BA",x"8C", -- 0x1158
		x"FC",x"D3",x"1D",x"57",x"8F",x"A1",x"C3",x"CD", -- 0x1160
		x"7B",x"9E",x"E3",x"57",x"F3",x"A4",x"05",x"10", -- 0x1168
		x"E1",x"FD",x"D6",x"71",x"0A",x"35",x"24",x"66", -- 0x1170
		x"80",x"97",x"E6",x"97",x"AD",x"21",x"A3",x"AA", -- 0x1178
		x"75",x"40",x"81",x"05",x"E2",x"C4",x"D2",x"DD", -- 0x1180
		x"64",x"36",x"35",x"D7",x"DA",x"3A",x"E8",x"BC", -- 0x1188
		x"B7",x"3F",x"AE",x"42",x"74",x"52",x"A8",x"F4", -- 0x1190
		x"E9",x"0F",x"0C",x"17",x"31",x"B0",x"42",x"A6", -- 0x1198
		x"F0",x"43",x"2B",x"D3",x"09",x"FD",x"32",x"EC", -- 0x11A0
		x"B4",x"67",x"C4",x"8F",x"22",x"2D",x"CC",x"D9", -- 0x11A8
		x"6D",x"FA",x"9B",x"E1",x"4D",x"45",x"57",x"37", -- 0x11B0
		x"54",x"63",x"CD",x"05",x"14",x"10",x"AB",x"85", -- 0x11B8
		x"54",x"D6",x"59",x"DC",x"55",x"0B",x"C9",x"0A", -- 0x11C0
		x"F2",x"0E",x"19",x"15",x"3C",x"65",x"6E",x"29", -- 0x11C8
		x"60",x"0B",x"0B",x"AD",x"50",x"E1",x"64",x"24", -- 0x11D0
		x"46",x"33",x"2A",x"5A",x"C2",x"55",x"DF",x"96", -- 0x11D8
		x"2D",x"B9",x"73",x"02",x"44",x"BC",x"8B",x"37", -- 0x11E0
		x"4B",x"24",x"4C",x"07",x"8A",x"3B",x"30",x"6A", -- 0x11E8
		x"46",x"BA",x"19",x"16",x"9D",x"7D",x"B9",x"E3", -- 0x11F0
		x"30",x"E3",x"BD",x"F3",x"3A",x"1E",x"8A",x"E6", -- 0x11F8
		x"57",x"7E",x"E8",x"9B",x"3B",x"F3",x"D3",x"86", -- 0x1200
		x"18",x"9F",x"0D",x"22",x"5A",x"3D",x"8D",x"A0", -- 0x1208
		x"78",x"A6",x"36",x"16",x"A3",x"F0",x"79",x"D4", -- 0x1210
		x"54",x"37",x"48",x"8E",x"D4",x"D2",x"F4",x"2C", -- 0x1218
		x"51",x"5D",x"C8",x"0D",x"51",x"1C",x"13",x"E9", -- 0x1220
		x"3B",x"21",x"0C",x"96",x"DD",x"99",x"B6",x"56", -- 0x1228
		x"BF",x"ED",x"EB",x"E3",x"5E",x"65",x"38",x"B2", -- 0x1230
		x"1D",x"80",x"C1",x"F1",x"D2",x"B6",x"9E",x"A4", -- 0x1238
		x"94",x"E6",x"B1",x"E5",x"03",x"44",x"4F",x"BD", -- 0x1240
		x"E4",x"DB",x"54",x"C3",x"75",x"0C",x"99",x"B5", -- 0x1248
		x"79",x"86",x"99",x"D7",x"6B",x"51",x"8A",x"08", -- 0x1250
		x"51",x"CB",x"FA",x"24",x"83",x"19",x"C8",x"18", -- 0x1258
		x"00",x"F9",x"7D",x"82",x"BE",x"4D",x"40",x"A3", -- 0x1260
		x"29",x"15",x"E6",x"1E",x"21",x"81",x"D3",x"1A", -- 0x1268
		x"87",x"EC",x"F1",x"F2",x"BD",x"FB",x"7B",x"0F", -- 0x1270
		x"C8",x"76",x"34",x"CB",x"0F",x"7C",x"63",x"0F", -- 0x1278
		x"F6",x"60",x"91",x"B5",x"AD",x"51",x"D8",x"D6", -- 0x1280
		x"66",x"C0",x"F5",x"07",x"C1",x"49",x"21",x"49", -- 0x1288
		x"B6",x"92",x"BB",x"74",x"8F",x"37",x"04",x"D7", -- 0x1290
		x"2D",x"38",x"23",x"3C",x"34",x"86",x"CA",x"2B", -- 0x1298
		x"E6",x"DB",x"60",x"95",x"2E",x"3A",x"EB",x"94", -- 0x12A0
		x"7A",x"61",x"9C",x"3C",x"2B",x"3D",x"05",x"E1", -- 0x12A8
		x"D0",x"C0",x"D5",x"DF",x"78",x"D9",x"B7",x"A5", -- 0x12B0
		x"91",x"DA",x"62",x"C6",x"61",x"2D",x"71",x"C7", -- 0x12B8
		x"0A",x"52",x"DC",x"38",x"0C",x"49",x"4C",x"86", -- 0x12C0
		x"AA",x"68",x"42",x"D5",x"A6",x"47",x"37",x"77", -- 0x12C8
		x"87",x"8D",x"57",x"00",x"E6",x"8E",x"A6",x"79", -- 0x12D0
		x"69",x"88",x"BF",x"4A",x"B5",x"B0",x"91",x"3F", -- 0x12D8
		x"03",x"6F",x"F6",x"0F",x"B8",x"44",x"15",x"E2", -- 0x12E0
		x"AC",x"57",x"39",x"53",x"1E",x"70",x"4A",x"A6", -- 0x12E8
		x"7D",x"21",x"A6",x"E4",x"AF",x"CC",x"DD",x"98", -- 0x12F0
		x"55",x"9D",x"E2",x"0C",x"CD",x"F4",x"4B",x"51", -- 0x12F8
		x"64",x"43",x"DF",x"9C",x"07",x"F5",x"7F",x"33", -- 0x1300
		x"CC",x"B8",x"07",x"EB",x"A9",x"51",x"92",x"A6", -- 0x1308
		x"73",x"B8",x"8B",x"A2",x"86",x"69",x"3C",x"DB", -- 0x1310
		x"86",x"9E",x"67",x"D4",x"93",x"33",x"26",x"77", -- 0x1318
		x"F5",x"06",x"14",x"FC",x"7B",x"14",x"30",x"49", -- 0x1320
		x"4C",x"37",x"B4",x"75",x"09",x"47",x"9C",x"7C", -- 0x1328
		x"00",x"A7",x"9E",x"86",x"91",x"DA",x"E2",x"18", -- 0x1330
		x"7A",x"4A",x"6C",x"0E",x"7D",x"92",x"06",x"F2", -- 0x1338
		x"19",x"99",x"EF",x"94",x"2D",x"A0",x"DD",x"7A", -- 0x1340
		x"D7",x"92",x"6F",x"60",x"59",x"8B",x"5C",x"D9", -- 0x1348
		x"34",x"FB",x"DF",x"C5",x"D6",x"C2",x"5D",x"D0", -- 0x1350
		x"8D",x"CA",x"DF",x"8A",x"DC",x"65",x"7E",x"F5", -- 0x1358
		x"FE",x"6E",x"8B",x"2D",x"0F",x"69",x"27",x"67", -- 0x1360
		x"7C",x"16",x"47",x"55",x"A2",x"A4",x"2F",x"D6", -- 0x1368
		x"A0",x"10",x"1C",x"F6",x"D2",x"79",x"C8",x"DF", -- 0x1370
		x"C3",x"28",x"6B",x"A1",x"8D",x"E9",x"97",x"0C", -- 0x1378
		x"58",x"23",x"39",x"E7",x"0D",x"DF",x"CE",x"09", -- 0x1380
		x"F6",x"95",x"5E",x"99",x"3A",x"8E",x"EF",x"5A", -- 0x1388
		x"9E",x"0C",x"52",x"F0",x"05",x"9A",x"D1",x"C9", -- 0x1390
		x"C2",x"3D",x"6B",x"CF",x"A6",x"82",x"DB",x"7E", -- 0x1398
		x"A6",x"95",x"E5",x"33",x"75",x"B4",x"3C",x"EB", -- 0x13A0
		x"4B",x"9A",x"05",x"05",x"A8",x"F4",x"60",x"C6", -- 0x13A8
		x"80",x"32",x"B8",x"06",x"4C",x"0A",x"4F",x"0F", -- 0x13B0
		x"C6",x"3A",x"5E",x"6D",x"BC",x"3A",x"EB",x"E2", -- 0x13B8
		x"4F",x"D2",x"16",x"45",x"07",x"D1",x"31",x"D1", -- 0x13C0
		x"EC",x"37",x"D7",x"95",x"AB",x"B7",x"5D",x"AC", -- 0x13C8
		x"69",x"95",x"B2",x"B5",x"9F",x"02",x"44",x"E5", -- 0x13D0
		x"3C",x"A2",x"53",x"78",x"5C",x"BE",x"5C",x"AC", -- 0x13D8
		x"91",x"F1",x"F1",x"19",x"44",x"23",x"EA",x"31", -- 0x13E0
		x"D9",x"42",x"46",x"86",x"F9",x"23",x"B2",x"E2", -- 0x13E8
		x"38",x"65",x"98",x"57",x"E6",x"DC",x"3D",x"A2", -- 0x13F0
		x"7F",x"10",x"1B",x"5C",x"CF",x"F6",x"09",x"61", -- 0x13F8
		x"69",x"7A",x"F9",x"AD",x"1D",x"E5",x"5E",x"F7", -- 0x1400
		x"28",x"24",x"FD",x"A2",x"48",x"B0",x"85",x"00", -- 0x1408
		x"95",x"9E",x"58",x"7C",x"7B",x"95",x"9E",x"7B", -- 0x1410
		x"26",x"39",x"D7",x"F5",x"B0",x"60",x"D6",x"1A", -- 0x1418
		x"DA",x"D1",x"C7",x"F7",x"B7",x"26",x"6F",x"5F", -- 0x1420
		x"4A",x"6D",x"81",x"12",x"9D",x"87",x"13",x"33", -- 0x1428
		x"26",x"EA",x"2F",x"21",x"00",x"4D",x"1C",x"26", -- 0x1430
		x"87",x"73",x"1C",x"38",x"D3",x"F3",x"52",x"2E", -- 0x1438
		x"C5",x"99",x"A6",x"FC",x"3F",x"16",x"DB",x"89", -- 0x1440
		x"04",x"DD",x"1C",x"A1",x"65",x"AE",x"55",x"0B", -- 0x1448
		x"99",x"84",x"2C",x"99",x"52",x"C8",x"C0",x"D9", -- 0x1450
		x"3C",x"5C",x"91",x"90",x"50",x"E3",x"3E",x"95", -- 0x1458
		x"FC",x"E4",x"12",x"3C",x"7B",x"6E",x"45",x"FE", -- 0x1460
		x"4C",x"61",x"20",x"B1",x"10",x"75",x"BC",x"29", -- 0x1468
		x"7A",x"68",x"C3",x"CC",x"B0",x"04",x"26",x"6D", -- 0x1470
		x"60",x"B7",x"FD",x"31",x"1B",x"BB",x"C6",x"18", -- 0x1478
		x"A1",x"59",x"D3",x"9C",x"C7",x"19",x"1B",x"14", -- 0x1480
		x"7B",x"3B",x"45",x"0B",x"31",x"81",x"35",x"2B", -- 0x1488
		x"69",x"78",x"77",x"1B",x"7C",x"1D",x"88",x"DC", -- 0x1490
		x"D4",x"06",x"8D",x"6F",x"C1",x"55",x"07",x"E2", -- 0x1498
		x"2E",x"DA",x"FE",x"F5",x"73",x"1A",x"89",x"6E", -- 0x14A0
		x"56",x"4E",x"7A",x"07",x"CF",x"2F",x"B1",x"B8", -- 0x14A8
		x"A7",x"29",x"D3",x"24",x"C5",x"DB",x"80",x"1A", -- 0x14B0
		x"61",x"0F",x"89",x"24",x"E3",x"10",x"86",x"12", -- 0x14B8
		x"6A",x"86",x"87",x"DD",x"A0",x"90",x"4D",x"76", -- 0x14C0
		x"DE",x"47",x"FC",x"2E",x"76",x"AE",x"E6",x"1E", -- 0x14C8
		x"57",x"BB",x"C1",x"1D",x"17",x"42",x"37",x"79", -- 0x14D0
		x"D0",x"40",x"1D",x"B4",x"CF",x"A3",x"46",x"3A", -- 0x14D8
		x"2A",x"4D",x"98",x"CB",x"DD",x"65",x"C1",x"3C", -- 0x14E0
		x"AC",x"BF",x"6A",x"A2",x"6E",x"52",x"C0",x"C6", -- 0x14E8
		x"8D",x"02",x"63",x"24",x"C3",x"9B",x"1D",x"95", -- 0x14F0
		x"5B",x"3A",x"C9",x"2C",x"DE",x"11",x"E5",x"88", -- 0x14F8
		x"DD",x"7E",x"D3",x"3C",x"E3",x"96",x"78",x"10", -- 0x1500
		x"56",x"63",x"B2",x"44",x"35",x"F2",x"0B",x"C2", -- 0x1508
		x"F4",x"EE",x"66",x"B9",x"0A",x"84",x"CE",x"65", -- 0x1510
		x"BE",x"98",x"91",x"1D",x"29",x"F7",x"A6",x"87", -- 0x1518
		x"76",x"7A",x"C3",x"DA",x"90",x"BB",x"EA",x"E6", -- 0x1520
		x"1F",x"9E",x"2C",x"54",x"11",x"B6",x"96",x"86", -- 0x1528
		x"A5",x"FD",x"BF",x"2F",x"02",x"8E",x"95",x"40", -- 0x1530
		x"A6",x"A6",x"5E",x"D0",x"9E",x"84",x"58",x"16", -- 0x1538
		x"7E",x"9B",x"F0",x"10",x"57",x"5B",x"76",x"77", -- 0x1540
		x"79",x"A2",x"4B",x"8B",x"D9",x"62",x"91",x"FE", -- 0x1548
		x"60",x"51",x"2F",x"E1",x"5F",x"44",x"22",x"06", -- 0x1550
		x"EA",x"00",x"56",x"0A",x"84",x"2E",x"20",x"83", -- 0x1558
		x"C9",x"90",x"93",x"22",x"6B",x"0A",x"19",x"E5", -- 0x1560
		x"2D",x"64",x"F0",x"86",x"46",x"82",x"85",x"A6", -- 0x1568
		x"53",x"34",x"08",x"B2",x"78",x"2B",x"B8",x"64", -- 0x1570
		x"AA",x"8F",x"6E",x"30",x"BD",x"0E",x"B3",x"08", -- 0x1578
		x"1E",x"C6",x"2A",x"09",x"50",x"C2",x"EE",x"FC", -- 0x1580
		x"A6",x"5F",x"83",x"ED",x"E1",x"89",x"14",x"35", -- 0x1588
		x"BD",x"1D",x"67",x"B6",x"C7",x"A0",x"9A",x"72", -- 0x1590
		x"30",x"88",x"22",x"6D",x"16",x"55",x"75",x"B3", -- 0x1598
		x"1C",x"1F",x"BC",x"EC",x"E1",x"2C",x"E9",x"89", -- 0x15A0
		x"8B",x"ED",x"F6",x"ED",x"77",x"0B",x"A2",x"B4", -- 0x15A8
		x"A7",x"0B",x"6B",x"EE",x"AB",x"85",x"62",x"5B", -- 0x15B0
		x"0E",x"04",x"C8",x"24",x"5A",x"3F",x"D7",x"F5", -- 0x15B8
		x"5E",x"95",x"E2",x"41",x"C1",x"CD",x"4A",x"4D", -- 0x15C0
		x"BB",x"C0",x"BA",x"B2",x"CB",x"5E",x"67",x"F3", -- 0x15C8
		x"69",x"53",x"E2",x"94",x"D8",x"C4",x"EF",x"E7", -- 0x15D0
		x"C9",x"38",x"8B",x"24",x"77",x"64",x"99",x"D6", -- 0x15D8
		x"79",x"7D",x"97",x"3B",x"CA",x"61",x"08",x"86", -- 0x15E0
		x"A1",x"C3",x"B8",x"EC",x"22",x"9F",x"E0",x"0B", -- 0x15E8
		x"72",x"44",x"1F",x"4C",x"09",x"0F",x"B3",x"52", -- 0x15F0
		x"47",x"BE",x"F5",x"3F",x"23",x"90",x"95",x"9C", -- 0x15F8
		x"0E",x"AC",x"57",x"D8",x"0E",x"60",x"DE",x"2F", -- 0x1600
		x"A3",x"97",x"1C",x"45",x"37",x"FD",x"50",x"AA", -- 0x1608
		x"42",x"6F",x"76",x"CA",x"FD",x"A9",x"1E",x"C4", -- 0x1610
		x"68",x"93",x"04",x"0C",x"24",x"99",x"A8",x"B1", -- 0x1618
		x"46",x"01",x"8A",x"D3",x"E0",x"E8",x"03",x"84", -- 0x1620
		x"80",x"20",x"C9",x"38",x"9D",x"99",x"62",x"5F", -- 0x1628
		x"88",x"58",x"2A",x"86",x"02",x"C7",x"4B",x"E9", -- 0x1630
		x"5C",x"CF",x"F5",x"00",x"69",x"1F",x"B2",x"30", -- 0x1638
		x"20",x"3D",x"83",x"80",x"A6",x"07",x"05",x"A6", -- 0x1640
		x"27",x"4E",x"DE",x"44",x"E7",x"C0",x"A3",x"70", -- 0x1648
		x"98",x"4D",x"76",x"1A",x"95",x"C1",x"05",x"71", -- 0x1650
		x"11",x"7A",x"71",x"7B",x"99",x"24",x"2B",x"39", -- 0x1658
		x"E1",x"AE",x"B9",x"88",x"B5",x"3E",x"2F",x"5C", -- 0x1660
		x"8C",x"8E",x"20",x"F3",x"CE",x"C3",x"E3",x"68", -- 0x1668
		x"91",x"5A",x"82",x"27",x"9C",x"87",x"98",x"AD", -- 0x1670
		x"03",x"89",x"A8",x"9C",x"AE",x"D3",x"56",x"90", -- 0x1678
		x"03",x"10",x"98",x"38",x"4F",x"47",x"95",x"5B", -- 0x1680
		x"D5",x"B5",x"CF",x"A5",x"F9",x"33",x"0E",x"0B", -- 0x1688
		x"0E",x"90",x"32",x"AA",x"98",x"4A",x"D7",x"1B", -- 0x1690
		x"D3",x"01",x"37",x"02",x"54",x"8D",x"12",x"57", -- 0x1698
		x"9E",x"AA",x"10",x"6D",x"F2",x"A5",x"48",x"48", -- 0x16A0
		x"DA",x"18",x"ED",x"54",x"4C",x"7B",x"5F",x"5A", -- 0x16A8
		x"8C",x"11",x"84",x"25",x"DA",x"DB",x"40",x"2F", -- 0x16B0
		x"5C",x"77",x"31",x"B1",x"06",x"44",x"88",x"24", -- 0x16B8
		x"6E",x"98",x"11",x"E0",x"BD",x"59",x"2A",x"19", -- 0x16C0
		x"F1",x"18",x"EC",x"BD",x"14",x"4D",x"97",x"A0", -- 0x16C8
		x"DD",x"1C",x"C5",x"39",x"77",x"85",x"68",x"D4", -- 0x16D0
		x"FC",x"19",x"06",x"82",x"5D",x"8E",x"A6",x"4C", -- 0x16D8
		x"A7",x"B7",x"2D",x"E4",x"91",x"57",x"FD",x"83", -- 0x16E0
		x"EF",x"EB",x"41",x"83",x"B8",x"D8",x"24",x"16", -- 0x16E8
		x"74",x"69",x"4F",x"6B",x"EE",x"37",x"40",x"6B", -- 0x16F0
		x"51",x"C5",x"EE",x"2E",x"D4",x"15",x"7A",x"7C", -- 0x16F8
		x"4D",x"28",x"E0",x"DE",x"FE",x"DF",x"E1",x"6E", -- 0x1700
		x"4B",x"23",x"F1",x"83",x"7B",x"16",x"19",x"EF", -- 0x1708
		x"7F",x"69",x"5B",x"6E",x"A0",x"1C",x"5A",x"71", -- 0x1710
		x"E1",x"49",x"A0",x"36",x"DD",x"9A",x"B2",x"2B", -- 0x1718
		x"C2",x"14",x"89",x"C2",x"73",x"6B",x"31",x"BE", -- 0x1720
		x"8E",x"24",x"C1",x"0A",x"B9",x"DA",x"79",x"B9", -- 0x1728
		x"C3",x"55",x"A7",x"65",x"71",x"02",x"56",x"D2", -- 0x1730
		x"4B",x"F6",x"0A",x"2A",x"92",x"3C",x"D4",x"D4", -- 0x1738
		x"50",x"5F",x"17",x"C3",x"4A",x"C8",x"02",x"59", -- 0x1740
		x"6C",x"C3",x"E2",x"26",x"1F",x"5D",x"DF",x"E2", -- 0x1748
		x"B2",x"88",x"C7",x"A3",x"8A",x"1F",x"76",x"56", -- 0x1750
		x"16",x"80",x"00",x"28",x"3D",x"54",x"7D",x"8D", -- 0x1758
		x"B3",x"94",x"D1",x"FE",x"5D",x"D3",x"D7",x"C9", -- 0x1760
		x"18",x"BA",x"70",x"37",x"18",x"50",x"1A",x"4A", -- 0x1768
		x"58",x"E2",x"ED",x"63",x"81",x"E4",x"B9",x"17", -- 0x1770
		x"65",x"39",x"40",x"22",x"8D",x"BD",x"B0",x"42", -- 0x1778
		x"D1",x"02",x"C0",x"30",x"D5",x"18",x"79",x"6D", -- 0x1780
		x"D2",x"E9",x"A4",x"EB",x"3B",x"3F",x"B5",x"13", -- 0x1788
		x"A1",x"A4",x"76",x"23",x"89",x"30",x"B9",x"6E", -- 0x1790
		x"69",x"F9",x"91",x"77",x"37",x"C1",x"39",x"89", -- 0x1798
		x"C3",x"79",x"B9",x"19",x"91",x"B2",x"87",x"64", -- 0x17A0
		x"9D",x"AB",x"CF",x"58",x"6A",x"86",x"6B",x"0C", -- 0x17A8
		x"2B",x"E2",x"AE",x"34",x"92",x"69",x"22",x"7C", -- 0x17B0
		x"E2",x"33",x"F3",x"9A",x"F4",x"2D",x"24",x"38", -- 0x17B8
		x"A6",x"5D",x"D1",x"38",x"10",x"59",x"9C",x"2D", -- 0x17C0
		x"84",x"6D",x"85",x"EF",x"73",x"F1",x"7B",x"9E", -- 0x17C8
		x"54",x"2B",x"52",x"E6",x"14",x"74",x"E2",x"76", -- 0x17D0
		x"28",x"D6",x"11",x"9C",x"83",x"B4",x"D5",x"2A", -- 0x17D8
		x"12",x"A7",x"E1",x"A2",x"80",x"FE",x"CF",x"84", -- 0x17E0
		x"EB",x"D5",x"74",x"5F",x"C7",x"70",x"7D",x"1C", -- 0x17E8
		x"1B",x"CF",x"82",x"2F",x"C3",x"66",x"A5",x"6B", -- 0x17F0
		x"BC",x"37",x"09",x"41",x"EB",x"DE",x"EA",x"7E", -- 0x17F8
		x"06",x"CD",x"A0",x"06",x"4C",x"EF",x"8A",x"38", -- 0x1800
		x"C5",x"7F",x"97",x"0D",x"6F",x"94",x"29",x"8A", -- 0x1808
		x"E3",x"2C",x"B9",x"A7",x"12",x"DE",x"93",x"CE", -- 0x1810
		x"16",x"9C",x"10",x"03",x"7B",x"FB",x"81",x"01", -- 0x1818
		x"49",x"22",x"86",x"95",x"91",x"90",x"4D",x"58", -- 0x1820
		x"10",x"64",x"65",x"7F",x"F8",x"0F",x"89",x"DC", -- 0x1828
		x"3B",x"43",x"04",x"4D",x"A2",x"97",x"9B",x"B8", -- 0x1830
		x"34",x"AC",x"BB",x"2F",x"28",x"BC",x"30",x"71", -- 0x1838
		x"5E",x"36",x"86",x"F0",x"C7",x"D3",x"49",x"57", -- 0x1840
		x"38",x"2E",x"57",x"B0",x"3D",x"E0",x"8D",x"F7", -- 0x1848
		x"A4",x"91",x"C4",x"47",x"2A",x"61",x"00",x"DD", -- 0x1850
		x"0E",x"3C",x"0E",x"36",x"F8",x"BD",x"27",x"D7", -- 0x1858
		x"F4",x"2D",x"48",x"3C",x"01",x"91",x"93",x"B8", -- 0x1860
		x"3F",x"EA",x"69",x"7D",x"CC",x"F6",x"75",x"71", -- 0x1868
		x"08",x"BA",x"B8",x"B1",x"1C",x"B8",x"90",x"A9", -- 0x1870
		x"74",x"1E",x"DF",x"6E",x"5B",x"86",x"C5",x"CF", -- 0x1878
		x"B3",x"0E",x"0C",x"34",x"1F",x"A0",x"6C",x"5E", -- 0x1880
		x"8B",x"55",x"5B",x"D7",x"4C",x"51",x"49",x"D3", -- 0x1888
		x"0C",x"81",x"06",x"28",x"BA",x"96",x"D1",x"2F", -- 0x1890
		x"34",x"31",x"1D",x"8F",x"37",x"E2",x"60",x"EA", -- 0x1898
		x"F0",x"EB",x"9E",x"8F",x"8C",x"8A",x"EE",x"98", -- 0x18A0
		x"DF",x"4A",x"70",x"AB",x"9B",x"BA",x"7F",x"A7", -- 0x18A8
		x"3C",x"85",x"4F",x"F6",x"9B",x"21",x"A6",x"CF", -- 0x18B0
		x"D1",x"C3",x"DF",x"09",x"A7",x"BF",x"73",x"18", -- 0x18B8
		x"AB",x"91",x"A8",x"B8",x"1C",x"17",x"51",x"FB", -- 0x18C0
		x"61",x"C1",x"A7",x"7D",x"FB",x"28",x"25",x"B8", -- 0x18C8
		x"2D",x"F4",x"2F",x"C9",x"16",x"D5",x"19",x"68", -- 0x18D0
		x"9A",x"78",x"71",x"C1",x"38",x"E5",x"D9",x"64", -- 0x18D8
		x"F6",x"02",x"1D",x"14",x"19",x"6E",x"10",x"FA", -- 0x18E0
		x"AF",x"B8",x"78",x"AC",x"60",x"1D",x"65",x"8D", -- 0x18E8
		x"12",x"94",x"D6",x"29",x"6B",x"70",x"11",x"85", -- 0x18F0
		x"68",x"82",x"47",x"A1",x"E7",x"A0",x"85",x"DF", -- 0x18F8
		x"23",x"A2",x"F3",x"3C",x"90",x"83",x"B6",x"40", -- 0x1900
		x"3C",x"2F",x"6C",x"1C",x"4D",x"51",x"2A",x"DE", -- 0x1908
		x"E6",x"80",x"87",x"D1",x"70",x"98",x"D6",x"D9", -- 0x1910
		x"1C",x"1E",x"FA",x"83",x"3E",x"80",x"63",x"61", -- 0x1918
		x"A2",x"D6",x"1E",x"B2",x"5B",x"D4",x"72",x"17", -- 0x1920
		x"84",x"DF",x"B3",x"51",x"31",x"DD",x"30",x"97", -- 0x1928
		x"5E",x"B8",x"69",x"CF",x"51",x"40",x"29",x"EC", -- 0x1930
		x"DD",x"24",x"71",x"9C",x"A4",x"D4",x"FD",x"C6", -- 0x1938
		x"2C",x"9B",x"79",x"87",x"F0",x"EB",x"1E",x"75", -- 0x1940
		x"4B",x"D1",x"46",x"FC",x"AF",x"76",x"94",x"8E", -- 0x1948
		x"AE",x"7E",x"DD",x"01",x"3E",x"07",x"ED",x"9C", -- 0x1950
		x"2B",x"5F",x"39",x"4F",x"B4",x"B6",x"16",x"E0", -- 0x1958
		x"53",x"0F",x"E7",x"44",x"7A",x"06",x"39",x"C6", -- 0x1960
		x"D8",x"7F",x"C3",x"08",x"75",x"D7",x"16",x"25", -- 0x1968
		x"56",x"F3",x"26",x"15",x"7A",x"93",x"B1",x"25", -- 0x1970
		x"73",x"EA",x"74",x"28",x"A1",x"0A",x"88",x"74", -- 0x1978
		x"98",x"70",x"38",x"14",x"76",x"F0",x"DA",x"CE", -- 0x1980
		x"EF",x"1E",x"57",x"66",x"F5",x"6D",x"8B",x"4D", -- 0x1988
		x"62",x"31",x"62",x"5C",x"44",x"93",x"82",x"B7", -- 0x1990
		x"7E",x"76",x"5F",x"9F",x"81",x"E7",x"94",x"1A", -- 0x1998
		x"58",x"CC",x"AD",x"4F",x"BE",x"88",x"1E",x"2E", -- 0x19A0
		x"26",x"75",x"94",x"1D",x"E3",x"9F",x"E9",x"C5", -- 0x19A8
		x"50",x"CB",x"22",x"95",x"5F",x"A4",x"CC",x"5D", -- 0x19B0
		x"1C",x"2D",x"FC",x"1D",x"94",x"91",x"B6",x"ED", -- 0x19B8
		x"DE",x"65",x"3D",x"1D",x"6D",x"DA",x"4B",x"14", -- 0x19C0
		x"D0",x"60",x"31",x"34",x"00",x"9A",x"F9",x"D0", -- 0x19C8
		x"66",x"9B",x"E5",x"C5",x"C0",x"B2",x"23",x"5C", -- 0x19D0
		x"5F",x"9F",x"F8",x"F4",x"B1",x"2F",x"62",x"90", -- 0x19D8
		x"14",x"1F",x"2D",x"82",x"79",x"78",x"16",x"4A", -- 0x19E0
		x"58",x"47",x"FD",x"59",x"E1",x"F7",x"2A",x"C7", -- 0x19E8
		x"14",x"8F",x"8D",x"54",x"42",x"30",x"30",x"22", -- 0x19F0
		x"CF",x"29",x"96",x"01",x"58",x"F8",x"11",x"6D", -- 0x19F8
		x"97",x"3E",x"6F",x"11",x"37",x"85",x"DB",x"8F", -- 0x1A00
		x"4C",x"D9",x"E8",x"AD",x"52",x"92",x"75",x"66", -- 0x1A08
		x"22",x"82",x"3A",x"E4",x"B2",x"6A",x"86",x"02", -- 0x1A10
		x"93",x"1D",x"83",x"6B",x"95",x"94",x"D8",x"2D", -- 0x1A18
		x"D3",x"C7",x"3E",x"0B",x"CC",x"99",x"1A",x"19", -- 0x1A20
		x"74",x"83",x"C6",x"C6",x"16",x"BB",x"AC",x"B8", -- 0x1A28
		x"3E",x"66",x"1D",x"70",x"D0",x"A3",x"F2",x"E3", -- 0x1A30
		x"40",x"76",x"4F",x"D5",x"0B",x"A8",x"03",x"5E", -- 0x1A38
		x"70",x"C0",x"69",x"3E",x"5B",x"84",x"D6",x"4F", -- 0x1A40
		x"08",x"1E",x"95",x"9D",x"D9",x"42",x"D5",x"98", -- 0x1A48
		x"A8",x"72",x"09",x"F8",x"16",x"7B",x"DC",x"56", -- 0x1A50
		x"F1",x"2C",x"AB",x"7D",x"54",x"AE",x"DB",x"45", -- 0x1A58
		x"EF",x"C5",x"03",x"CA",x"4A",x"D9",x"1A",x"D1", -- 0x1A60
		x"F7",x"AF",x"EE",x"52",x"71",x"C5",x"EA",x"99", -- 0x1A68
		x"B7",x"73",x"92",x"CE",x"6F",x"EE",x"A4",x"E0", -- 0x1A70
		x"9A",x"D0",x"5E",x"EF",x"FE",x"BA",x"35",x"EE", -- 0x1A78
		x"80",x"38",x"39",x"4A",x"91",x"D2",x"1C",x"0A", -- 0x1A80
		x"02",x"8A",x"5C",x"F2",x"CF",x"C6",x"8C",x"88", -- 0x1A88
		x"B9",x"9E",x"D6",x"29",x"8D",x"FA",x"0B",x"29", -- 0x1A90
		x"CB",x"E8",x"19",x"CB",x"A3",x"CD",x"3A",x"24", -- 0x1A98
		x"85",x"F3",x"6E",x"17",x"C6",x"0A",x"21",x"C9", -- 0x1AA0
		x"95",x"FC",x"BC",x"E4",x"C3",x"C9",x"6D",x"7E", -- 0x1AA8
		x"68",x"C3",x"27",x"76",x"BF",x"32",x"9F",x"0B", -- 0x1AB0
		x"1C",x"38",x"56",x"BF",x"85",x"91",x"64",x"0B", -- 0x1AB8
		x"05",x"D2",x"A1",x"CB",x"5D",x"43",x"15",x"72", -- 0x1AC0
		x"40",x"52",x"57",x"84",x"1C",x"45",x"82",x"04", -- 0x1AC8
		x"88",x"A9",x"7A",x"C7",x"5C",x"1A",x"D3",x"F7", -- 0x1AD0
		x"D1",x"2A",x"37",x"57",x"3B",x"9B",x"E1",x"40", -- 0x1AD8
		x"EE",x"84",x"8C",x"4C",x"47",x"A1",x"BE",x"87", -- 0x1AE0
		x"F3",x"95",x"8B",x"8F",x"5A",x"0E",x"94",x"E3", -- 0x1AE8
		x"38",x"0F",x"AB",x"94",x"A9",x"FE",x"0C",x"7B", -- 0x1AF0
		x"A9",x"43",x"53",x"64",x"5F",x"35",x"25",x"4E", -- 0x1AF8
		x"39",x"B1",x"1A",x"00",x"D2",x"58",x"08",x"C7", -- 0x1B00
		x"ED",x"93",x"57",x"C8",x"22",x"EB",x"AC",x"5A", -- 0x1B08
		x"7B",x"D7",x"6E",x"25",x"D7",x"F9",x"A0",x"81", -- 0x1B10
		x"3D",x"73",x"E5",x"9C",x"29",x"0B",x"6A",x"E1", -- 0x1B18
		x"3C",x"84",x"E2",x"10",x"DC",x"EA",x"57",x"4B", -- 0x1B20
		x"FD",x"AE",x"14",x"20",x"1B",x"40",x"F9",x"96", -- 0x1B28
		x"18",x"E7",x"3B",x"EF",x"E1",x"5B",x"F0",x"9F", -- 0x1B30
		x"CF",x"57",x"BB",x"F8",x"62",x"27",x"DA",x"1F", -- 0x1B38
		x"2B",x"3D",x"2F",x"88",x"28",x"86",x"D3",x"27", -- 0x1B40
		x"B4",x"67",x"C6",x"4F",x"A7",x"C1",x"65",x"BF", -- 0x1B48
		x"29",x"A0",x"30",x"0C",x"FC",x"21",x"AB",x"CC", -- 0x1B50
		x"78",x"E6",x"45",x"5B",x"0E",x"9F",x"7A",x"3A", -- 0x1B58
		x"DD",x"29",x"C2",x"85",x"2F",x"16",x"2C",x"E3", -- 0x1B60
		x"7D",x"F3",x"34",x"25",x"35",x"99",x"64",x"5E", -- 0x1B68
		x"BA",x"94",x"E9",x"B7",x"36",x"15",x"84",x"2E", -- 0x1B70
		x"FC",x"49",x"89",x"0B",x"E8",x"83",x"C4",x"46", -- 0x1B78
		x"2C",x"07",x"CC",x"5B",x"9C",x"F8",x"40",x"1A", -- 0x1B80
		x"EC",x"F3",x"BE",x"A1",x"0D",x"A3",x"01",x"C7", -- 0x1B88
		x"38",x"EA",x"FE",x"ED",x"80",x"03",x"1D",x"7D", -- 0x1B90
		x"4C",x"26",x"08",x"B5",x"2A",x"4D",x"FB",x"56", -- 0x1B98
		x"D3",x"C8",x"B2",x"71",x"C2",x"72",x"0B",x"2F", -- 0x1BA0
		x"E5",x"4A",x"D1",x"72",x"ED",x"52",x"BA",x"A5", -- 0x1BA8
		x"BC",x"B9",x"94",x"3D",x"BD",x"B1",x"BA",x"0A", -- 0x1BB0
		x"57",x"43",x"BF",x"81",x"90",x"3C",x"D8",x"64", -- 0x1BB8
		x"05",x"0B",x"55",x"47",x"FC",x"61",x"77",x"E2", -- 0x1BC0
		x"2B",x"C8",x"55",x"19",x"1B",x"8F",x"BE",x"D7", -- 0x1BC8
		x"4A",x"D2",x"95",x"08",x"04",x"CF",x"91",x"5C", -- 0x1BD0
		x"13",x"D1",x"5D",x"A3",x"0E",x"36",x"88",x"13", -- 0x1BD8
		x"C0",x"DD",x"5B",x"BD",x"BE",x"52",x"20",x"E9", -- 0x1BE0
		x"1B",x"F5",x"82",x"36",x"85",x"C1",x"8D",x"CF", -- 0x1BE8
		x"94",x"23",x"57",x"19",x"F3",x"E9",x"75",x"86", -- 0x1BF0
		x"BB",x"D2",x"AA",x"C9",x"89",x"33",x"5C",x"C9", -- 0x1BF8
		x"90",x"37",x"88",x"CF",x"89",x"28",x"39",x"24", -- 0x1C00
		x"1E",x"BC",x"D9",x"A4",x"7E",x"68",x"F3",x"92", -- 0x1C08
		x"0B",x"4C",x"AB",x"FE",x"36",x"A0",x"06",x"71", -- 0x1C10
		x"F3",x"B0",x"BA",x"7D",x"E3",x"17",x"C6",x"F3", -- 0x1C18
		x"CE",x"4F",x"C3",x"58",x"78",x"FD",x"7D",x"16", -- 0x1C20
		x"3A",x"57",x"BA",x"B8",x"3F",x"AF",x"CA",x"4B", -- 0x1C28
		x"7B",x"77",x"C9",x"B1",x"97",x"CF",x"A2",x"8B", -- 0x1C30
		x"80",x"5D",x"88",x"E3",x"F3",x"50",x"D8",x"C2", -- 0x1C38
		x"1F",x"1C",x"1C",x"97",x"99",x"19",x"2E",x"D3", -- 0x1C40
		x"EF",x"E8",x"0C",x"30",x"18",x"D7",x"FA",x"13", -- 0x1C48
		x"CE",x"C4",x"44",x"66",x"15",x"E6",x"F2",x"95", -- 0x1C50
		x"C3",x"7B",x"F9",x"B8",x"4B",x"D2",x"7B",x"6B", -- 0x1C58
		x"6E",x"17",x"82",x"09",x"AF",x"B0",x"DC",x"A0", -- 0x1C60
		x"1A",x"69",x"50",x"32",x"C0",x"4B",x"C5",x"8F", -- 0x1C68
		x"8F",x"0A",x"75",x"A4",x"F1",x"68",x"BA",x"B5", -- 0x1C70
		x"64",x"B4",x"6E",x"2F",x"07",x"6A",x"9A",x"F4", -- 0x1C78
		x"01",x"1E",x"FD",x"B1",x"CE",x"5B",x"D1",x"68", -- 0x1C80
		x"C4",x"22",x"1B",x"85",x"EC",x"E0",x"94",x"7C", -- 0x1C88
		x"EA",x"0A",x"A1",x"DC",x"F2",x"DB",x"13",x"57", -- 0x1C90
		x"10",x"01",x"86",x"96",x"6B",x"A1",x"8B",x"6D", -- 0x1C98
		x"BF",x"8A",x"9E",x"0E",x"65",x"70",x"F6",x"2A", -- 0x1CA0
		x"92",x"12",x"2F",x"FE",x"F2",x"C3",x"FA",x"DD", -- 0x1CA8
		x"CD",x"9C",x"3B",x"C0",x"F7",x"CD",x"97",x"87", -- 0x1CB0
		x"CE",x"9E",x"1E",x"BA",x"BF",x"AA",x"A7",x"FE", -- 0x1CB8
		x"B4",x"46",x"0D",x"1A",x"B6",x"04",x"C3",x"C8", -- 0x1CC0
		x"95",x"F2",x"C7",x"88",x"36",x"C2",x"E6",x"04", -- 0x1CC8
		x"DF",x"22",x"45",x"D7",x"EF",x"5C",x"60",x"BE", -- 0x1CD0
		x"7A",x"FD",x"F8",x"3A",x"28",x"A0",x"39",x"DC", -- 0x1CD8
		x"E6",x"C6",x"76",x"9D",x"4A",x"B9",x"E5",x"E0", -- 0x1CE0
		x"AC",x"AD",x"69",x"62",x"71",x"CF",x"E6",x"51", -- 0x1CE8
		x"F1",x"2C",x"A8",x"61",x"08",x"88",x"A0",x"83", -- 0x1CF0
		x"07",x"99",x"3D",x"2F",x"3B",x"F6",x"8C",x"22", -- 0x1CF8
		x"BD",x"03",x"40",x"87",x"BD",x"26",x"68",x"E9", -- 0x1D00
		x"54",x"52",x"4D",x"C5",x"22",x"34",x"96",x"94", -- 0x1D08
		x"DF",x"BE",x"F5",x"67",x"C7",x"16",x"6A",x"CE", -- 0x1D10
		x"B0",x"A8",x"FD",x"EB",x"1F",x"0A",x"8D",x"DC", -- 0x1D18
		x"8D",x"4D",x"64",x"CA",x"F3",x"4D",x"B4",x"48", -- 0x1D20
		x"1F",x"81",x"8D",x"C0",x"35",x"24",x"55",x"94", -- 0x1D28
		x"62",x"CB",x"FC",x"2A",x"E1",x"E6",x"F8",x"92", -- 0x1D30
		x"0F",x"77",x"FD",x"2E",x"81",x"0C",x"0B",x"0F", -- 0x1D38
		x"D8",x"EF",x"D9",x"CC",x"BC",x"0F",x"15",x"DB", -- 0x1D40
		x"10",x"A2",x"9C",x"C5",x"46",x"72",x"5A",x"A9", -- 0x1D48
		x"3E",x"D6",x"D3",x"20",x"BE",x"4D",x"33",x"4D", -- 0x1D50
		x"44",x"31",x"7C",x"C5",x"BC",x"07",x"55",x"96", -- 0x1D58
		x"F6",x"AE",x"63",x"33",x"3D",x"F8",x"0F",x"4E", -- 0x1D60
		x"1B",x"2C",x"93",x"62",x"9E",x"ED",x"8B",x"DC", -- 0x1D68
		x"45",x"DE",x"7C",x"83",x"2C",x"AF",x"D0",x"70", -- 0x1D70
		x"61",x"4D",x"B6",x"9D",x"55",x"8B",x"34",x"CB", -- 0x1D78
		x"B9",x"18",x"00",x"F7",x"90",x"8E",x"C5",x"AB", -- 0x1D80
		x"3A",x"59",x"8D",x"D8",x"C6",x"19",x"35",x"8B", -- 0x1D88
		x"F8",x"B2",x"0F",x"A4",x"E1",x"E0",x"95",x"43", -- 0x1D90
		x"2E",x"CB",x"E1",x"03",x"57",x"95",x"4F",x"90", -- 0x1D98
		x"2D",x"CE",x"08",x"BD",x"5D",x"4D",x"6A",x"18", -- 0x1DA0
		x"26",x"F7",x"F0",x"ED",x"91",x"A6",x"79",x"8A", -- 0x1DA8
		x"59",x"89",x"AE",x"BA",x"E9",x"44",x"FE",x"97", -- 0x1DB0
		x"10",x"60",x"9B",x"E6",x"75",x"EA",x"F7",x"A3", -- 0x1DB8
		x"B9",x"00",x"61",x"96",x"4E",x"4B",x"AE",x"74", -- 0x1DC0
		x"C3",x"20",x"E1",x"55",x"C6",x"DB",x"5F",x"9F", -- 0x1DC8
		x"65",x"8D",x"5A",x"CE",x"D2",x"D8",x"66",x"62", -- 0x1DD0
		x"B8",x"81",x"C9",x"2F",x"6C",x"C1",x"52",x"A5", -- 0x1DD8
		x"C1",x"33",x"BC",x"8F",x"FE",x"EA",x"05",x"C2", -- 0x1DE0
		x"8A",x"E6",x"97",x"51",x"C2",x"76",x"70",x"A7", -- 0x1DE8
		x"04",x"CB",x"76",x"56",x"A4",x"5D",x"39",x"DD", -- 0x1DF0
		x"DE",x"03",x"8C",x"CB",x"44",x"DE",x"F0",x"06", -- 0x1DF8
		x"91",x"AD",x"96",x"90",x"19",x"1B",x"D2",x"A3", -- 0x1E00
		x"81",x"6A",x"75",x"45",x"60",x"E5",x"6C",x"65", -- 0x1E08
		x"31",x"63",x"3B",x"56",x"C0",x"74",x"34",x"9F", -- 0x1E10
		x"F6",x"C0",x"EA",x"3B",x"1F",x"DC",x"C1",x"30", -- 0x1E18
		x"0A",x"D7",x"C1",x"23",x"F2",x"14",x"47",x"74", -- 0x1E20
		x"FE",x"BC",x"39",x"5F",x"22",x"A6",x"44",x"D3", -- 0x1E28
		x"89",x"00",x"2A",x"4A",x"74",x"DD",x"69",x"6C", -- 0x1E30
		x"1E",x"D4",x"27",x"BC",x"B1",x"E8",x"EC",x"BB", -- 0x1E38
		x"C0",x"2E",x"5F",x"33",x"43",x"A6",x"28",x"C1", -- 0x1E40
		x"E2",x"61",x"21",x"05",x"87",x"E5",x"58",x"90", -- 0x1E48
		x"E5",x"82",x"DA",x"D9",x"60",x"C4",x"C5",x"FD", -- 0x1E50
		x"99",x"ED",x"BA",x"CA",x"56",x"A8",x"86",x"97", -- 0x1E58
		x"56",x"E5",x"CA",x"99",x"8C",x"72",x"5B",x"EE", -- 0x1E60
		x"54",x"FC",x"74",x"DB",x"62",x"CC",x"6D",x"48", -- 0x1E68
		x"50",x"C7",x"22",x"30",x"0C",x"68",x"2F",x"25", -- 0x1E70
		x"56",x"69",x"EF",x"AC",x"12",x"77",x"44",x"69", -- 0x1E78
		x"DC",x"8F",x"82",x"E9",x"02",x"5E",x"D8",x"56", -- 0x1E80
		x"DA",x"4D",x"B2",x"3D",x"1B",x"9F",x"05",x"EA", -- 0x1E88
		x"67",x"A6",x"9A",x"F3",x"0F",x"49",x"19",x"E4", -- 0x1E90
		x"B3",x"0A",x"92",x"C5",x"01",x"56",x"AE",x"5D", -- 0x1E98
		x"65",x"B1",x"47",x"68",x"8F",x"A0",x"3E",x"6A", -- 0x1EA0
		x"ED",x"70",x"27",x"88",x"10",x"2C",x"73",x"F7", -- 0x1EA8
		x"52",x"0F",x"EB",x"62",x"58",x"84",x"47",x"8B", -- 0x1EB0
		x"8E",x"59",x"D1",x"0F",x"30",x"80",x"6D",x"95", -- 0x1EB8
		x"B1",x"34",x"7D",x"41",x"D4",x"BC",x"2B",x"43", -- 0x1EC0
		x"AC",x"52",x"CB",x"BD",x"FD",x"BF",x"B5",x"51", -- 0x1EC8
		x"CE",x"21",x"33",x"A6",x"A5",x"F9",x"33",x"B4", -- 0x1ED0
		x"54",x"05",x"43",x"04",x"05",x"30",x"99",x"B7", -- 0x1ED8
		x"65",x"97",x"78",x"3A",x"D3",x"A4",x"7D",x"80", -- 0x1EE0
		x"F6",x"C9",x"3E",x"F5",x"89",x"73",x"C6",x"58", -- 0x1EE8
		x"94",x"F9",x"7E",x"BA",x"F3",x"31",x"6F",x"C7", -- 0x1EF0
		x"B5",x"32",x"CB",x"3B",x"63",x"E5",x"72",x"C8", -- 0x1EF8
		x"7D",x"EA",x"82",x"51",x"8F",x"80",x"D1",x"07", -- 0x1F00
		x"4A",x"11",x"7C",x"D3",x"04",x"43",x"AB",x"19", -- 0x1F08
		x"BC",x"A9",x"D3",x"B0",x"5B",x"C2",x"79",x"11", -- 0x1F10
		x"F4",x"C4",x"4C",x"58",x"AA",x"3E",x"A0",x"28", -- 0x1F18
		x"2A",x"24",x"79",x"39",x"24",x"CB",x"BF",x"6E", -- 0x1F20
		x"5C",x"3C",x"C1",x"60",x"FE",x"6D",x"79",x"BB", -- 0x1F28
		x"96",x"4D",x"EC",x"F1",x"8F",x"66",x"04",x"85", -- 0x1F30
		x"AA",x"CF",x"5D",x"56",x"0F",x"7E",x"7E",x"B8", -- 0x1F38
		x"22",x"78",x"F1",x"46",x"44",x"32",x"34",x"A0", -- 0x1F40
		x"ED",x"F5",x"80",x"ED",x"E2",x"FA",x"29",x"79", -- 0x1F48
		x"C7",x"16",x"6C",x"D7",x"FB",x"70",x"DC",x"A7", -- 0x1F50
		x"BF",x"3A",x"FD",x"4E",x"38",x"FB",x"07",x"5A", -- 0x1F58
		x"F3",x"79",x"A0",x"B7",x"AB",x"D4",x"D7",x"99", -- 0x1F60
		x"4A",x"59",x"07",x"2D",x"D3",x"31",x"A7",x"1B", -- 0x1F68
		x"47",x"14",x"F2",x"C3",x"04",x"CF",x"6B",x"C3", -- 0x1F70
		x"8A",x"E8",x"92",x"C2",x"64",x"99",x"9D",x"59", -- 0x1F78
		x"92",x"3E",x"11",x"3E",x"93",x"E9",x"58",x"DD", -- 0x1F80
		x"C2",x"5F",x"0C",x"96",x"10",x"B3",x"31",x"D7", -- 0x1F88
		x"C7",x"25",x"9B",x"4B",x"74",x"86",x"8E",x"7E", -- 0x1F90
		x"6F",x"21",x"C1",x"D3",x"BB",x"5F",x"AC",x"4E", -- 0x1F98
		x"1D",x"3E",x"0D",x"B0",x"28",x"E4",x"0F",x"6A", -- 0x1FA0
		x"44",x"1B",x"01",x"D4",x"4E",x"B1",x"AC",x"95", -- 0x1FA8
		x"D6",x"48",x"E0",x"CB",x"4E",x"6F",x"C9",x"BD", -- 0x1FB0
		x"91",x"8B",x"11",x"CC",x"EA",x"3E",x"9A",x"88", -- 0x1FB8
		x"7C",x"A7",x"39",x"24",x"0C",x"48",x"8E",x"D0", -- 0x1FC0
		x"E2",x"0F",x"A5",x"31",x"C0",x"52",x"C6",x"18", -- 0x1FC8
		x"1A",x"A7",x"63",x"68",x"97",x"2D",x"A5",x"A8", -- 0x1FD0
		x"B9",x"36",x"75",x"24",x"74",x"10",x"AC",x"70", -- 0x1FD8
		x"38",x"66",x"14",x"44",x"AE",x"A2",x"94",x"12", -- 0x1FE0
		x"31",x"3A",x"43",x"F2",x"0C",x"0B",x"8A",x"A5", -- 0x1FE8
		x"32",x"ED",x"8D",x"C9",x"1B",x"B2",x"F1",x"54", -- 0x1FF0
		x"E9",x"67",x"79",x"DD",x"F7",x"A5",x"CE",x"AF", -- 0x1FF8
		x"0C",x"E2",x"73",x"3B",x"86",x"09",x"4D",x"37", -- 0x2000
		x"43",x"10",x"2A",x"CF",x"9A",x"34",x"75",x"CD", -- 0x2008
		x"22",x"04",x"17",x"3E",x"36",x"0A",x"12",x"20", -- 0x2010
		x"F0",x"8B",x"7E",x"E8",x"B1",x"4D",x"98",x"3D", -- 0x2018
		x"30",x"8C",x"F7",x"36",x"95",x"C4",x"ED",x"58", -- 0x2020
		x"D5",x"97",x"28",x"70",x"CC",x"9E",x"BD",x"EE", -- 0x2028
		x"22",x"55",x"AC",x"58",x"DE",x"BF",x"F8",x"CF", -- 0x2030
		x"CA",x"F6",x"39",x"7C",x"44",x"51",x"3A",x"F3", -- 0x2038
		x"DD",x"32",x"AA",x"73",x"F7",x"98",x"CC",x"4D", -- 0x2040
		x"30",x"74",x"BD",x"FC",x"92",x"FB",x"6C",x"34", -- 0x2048
		x"51",x"19",x"0D",x"AF",x"58",x"06",x"7F",x"24", -- 0x2050
		x"FC",x"38",x"20",x"C0",x"8A",x"D9",x"B4",x"E7", -- 0x2058
		x"0D",x"DE",x"DB",x"84",x"77",x"A8",x"D1",x"28", -- 0x2060
		x"9C",x"8F",x"25",x"30",x"0B",x"11",x"64",x"DB", -- 0x2068
		x"2B",x"71",x"8B",x"03",x"F6",x"0C",x"A6",x"F3", -- 0x2070
		x"C3",x"C7",x"B4",x"4E",x"21",x"E9",x"B6",x"2E", -- 0x2078
		x"C8",x"92",x"B2",x"C0",x"BA",x"84",x"E8",x"57", -- 0x2080
		x"94",x"8D",x"87",x"9F",x"9F",x"6C",x"FB",x"4A", -- 0x2088
		x"DD",x"87",x"4D",x"55",x"13",x"F4",x"49",x"D7", -- 0x2090
		x"3C",x"7E",x"A5",x"5D",x"E7",x"5C",x"0C",x"30", -- 0x2098
		x"EE",x"BE",x"70",x"29",x"C3",x"59",x"81",x"D7", -- 0x20A0
		x"67",x"88",x"F6",x"07",x"F4",x"F2",x"D0",x"53", -- 0x20A8
		x"7B",x"9D",x"A8",x"8E",x"92",x"71",x"E5",x"4E", -- 0x20B0
		x"6F",x"8C",x"2C",x"57",x"68",x"38",x"08",x"D7", -- 0x20B8
		x"76",x"78",x"01",x"B9",x"D2",x"02",x"91",x"3A", -- 0x20C0
		x"8B",x"89",x"C0",x"00",x"FB",x"11",x"53",x"77", -- 0x20C8
		x"AE",x"7B",x"86",x"42",x"ED",x"6C",x"10",x"5D", -- 0x20D0
		x"78",x"3C",x"35",x"61",x"F3",x"3D",x"B8",x"EA", -- 0x20D8
		x"B5",x"B9",x"A4",x"08",x"3C",x"B6",x"C1",x"C7", -- 0x20E0
		x"40",x"02",x"47",x"3C",x"13",x"1B",x"34",x"C2", -- 0x20E8
		x"96",x"BA",x"84",x"04",x"A6",x"94",x"E1",x"9F", -- 0x20F0
		x"51",x"17",x"80",x"C4",x"D3",x"39",x"AF",x"89", -- 0x20F8
		x"72",x"D4",x"12",x"AE",x"8B",x"D3",x"F5",x"4B", -- 0x2100
		x"56",x"3E",x"07",x"69",x"59",x"3B",x"2C",x"6F", -- 0x2108
		x"75",x"30",x"74",x"9C",x"45",x"56",x"BB",x"96", -- 0x2110
		x"6D",x"3C",x"DA",x"C0",x"F4",x"0B",x"4A",x"E6", -- 0x2118
		x"5F",x"DB",x"96",x"EA",x"30",x"0C",x"B5",x"86", -- 0x2120
		x"C9",x"BC",x"EF",x"A2",x"F8",x"9C",x"13",x"ED", -- 0x2128
		x"CC",x"07",x"0A",x"12",x"5D",x"C5",x"28",x"4A", -- 0x2130
		x"81",x"83",x"0B",x"F5",x"8E",x"D4",x"DD",x"ED", -- 0x2138
		x"B1",x"F3",x"58",x"E1",x"7F",x"0E",x"E7",x"4A", -- 0x2140
		x"CA",x"D7",x"EC",x"43",x"F3",x"7F",x"B1",x"41", -- 0x2148
		x"86",x"BB",x"53",x"E3",x"02",x"FB",x"AD",x"83", -- 0x2150
		x"7F",x"B8",x"F9",x"8D",x"0E",x"D7",x"7B",x"3F", -- 0x2158
		x"4B",x"D3",x"A0",x"CA",x"61",x"88",x"15",x"AB", -- 0x2160
		x"DF",x"82",x"EF",x"D4",x"02",x"21",x"16",x"09", -- 0x2168
		x"DC",x"E8",x"EC",x"DE",x"E4",x"1B",x"E2",x"E3", -- 0x2170
		x"53",x"5C",x"71",x"61",x"34",x"6C",x"20",x"7F", -- 0x2178
		x"40",x"C0",x"4A",x"21",x"C8",x"DF",x"CD",x"A9", -- 0x2180
		x"62",x"BD",x"FD",x"E3",x"5E",x"93",x"EC",x"3B", -- 0x2188
		x"FB",x"5A",x"9A",x"61",x"75",x"FC",x"45",x"48", -- 0x2190
		x"59",x"B7",x"AA",x"0D",x"24",x"4A",x"0C",x"E4", -- 0x2198
		x"8B",x"56",x"85",x"54",x"B5",x"53",x"7D",x"18", -- 0x21A0
		x"90",x"FA",x"7C",x"EE",x"8E",x"69",x"AA",x"0B", -- 0x21A8
		x"C3",x"45",x"6C",x"B8",x"C1",x"B1",x"02",x"1B", -- 0x21B0
		x"E8",x"2C",x"28",x"8D",x"F5",x"B3",x"F1",x"81", -- 0x21B8
		x"0A",x"77",x"D6",x"40",x"4B",x"D3",x"58",x"DB", -- 0x21C0
		x"CF",x"54",x"CB",x"DD",x"BE",x"76",x"E8",x"02", -- 0x21C8
		x"3B",x"55",x"3B",x"FC",x"87",x"BC",x"97",x"70", -- 0x21D0
		x"E8",x"3F",x"7D",x"DE",x"F2",x"EE",x"E0",x"7C", -- 0x21D8
		x"67",x"B7",x"BC",x"B2",x"8B",x"95",x"0E",x"5B", -- 0x21E0
		x"E9",x"59",x"3A",x"28",x"4F",x"A2",x"AA",x"8A", -- 0x21E8
		x"F8",x"E5",x"07",x"80",x"A2",x"9E",x"70",x"0B", -- 0x21F0
		x"5D",x"6E",x"69",x"50",x"5D",x"4A",x"4D",x"44", -- 0x21F8
		x"02",x"0A",x"76",x"0E",x"1F",x"85",x"E8",x"89", -- 0x2200
		x"DE",x"A2",x"B1",x"AE",x"46",x"5C",x"B8",x"3F", -- 0x2208
		x"42",x"C0",x"3F",x"64",x"DE",x"AF",x"6F",x"3D", -- 0x2210
		x"1E",x"D9",x"0D",x"7C",x"A3",x"5A",x"40",x"A6", -- 0x2218
		x"E4",x"B7",x"34",x"04",x"3D",x"9C",x"8D",x"9B", -- 0x2220
		x"40",x"BF",x"4A",x"86",x"1C",x"04",x"45",x"DE", -- 0x2228
		x"44",x"84",x"43",x"23",x"B3",x"33",x"DF",x"52", -- 0x2230
		x"0D",x"6D",x"4E",x"B0",x"C7",x"8E",x"D6",x"2C", -- 0x2238
		x"46",x"8A",x"B0",x"03",x"28",x"BD",x"9F",x"68", -- 0x2240
		x"7D",x"69",x"6E",x"1A",x"EC",x"33",x"F8",x"31", -- 0x2248
		x"37",x"BB",x"D4",x"6A",x"EE",x"34",x"BC",x"7B", -- 0x2250
		x"A1",x"8A",x"AC",x"E9",x"1A",x"03",x"16",x"DF", -- 0x2258
		x"8E",x"46",x"E3",x"36",x"05",x"03",x"1E",x"82", -- 0x2260
		x"EB",x"8C",x"1C",x"D9",x"3F",x"15",x"8A",x"76", -- 0x2268
		x"D1",x"5F",x"E0",x"40",x"94",x"1E",x"BC",x"B5", -- 0x2270
		x"A8",x"69",x"9F",x"42",x"6C",x"36",x"23",x"7A", -- 0x2278
		x"7C",x"86",x"B0",x"81",x"89",x"CE",x"84",x"F4", -- 0x2280
		x"DA",x"A0",x"CE",x"1A",x"36",x"D9",x"10",x"87", -- 0x2288
		x"B8",x"71",x"C7",x"CC",x"8F",x"04",x"83",x"B7", -- 0x2290
		x"EC",x"23",x"FA",x"5A",x"59",x"1E",x"54",x"D6", -- 0x2298
		x"24",x"06",x"D7",x"AD",x"54",x"5C",x"22",x"AF", -- 0x22A0
		x"7D",x"71",x"C9",x"B3",x"4B",x"5A",x"BA",x"04", -- 0x22A8
		x"CB",x"82",x"D1",x"DA",x"07",x"55",x"92",x"F3", -- 0x22B0
		x"F7",x"8D",x"CD",x"52",x"2B",x"23",x"A8",x"4F", -- 0x22B8
		x"A8",x"80",x"7C",x"FC",x"DD",x"9F",x"AC",x"DA", -- 0x22C0
		x"11",x"F6",x"8E",x"DB",x"51",x"49",x"DF",x"9C", -- 0x22C8
		x"4B",x"31",x"77",x"52",x"06",x"0A",x"C6",x"FE", -- 0x22D0
		x"98",x"94",x"D0",x"43",x"B7",x"79",x"93",x"DF", -- 0x22D8
		x"F9",x"8F",x"5D",x"57",x"2F",x"89",x"32",x"BF", -- 0x22E0
		x"80",x"40",x"9B",x"51",x"09",x"FB",x"ED",x"D4", -- 0x22E8
		x"AC",x"E4",x"A6",x"B3",x"EF",x"6D",x"32",x"08", -- 0x22F0
		x"03",x"03",x"4B",x"3A",x"7C",x"5E",x"1B",x"F5", -- 0x22F8
		x"6E",x"78",x"4E",x"1D",x"81",x"00",x"DD",x"03", -- 0x2300
		x"C0",x"F8",x"D3",x"C9",x"74",x"42",x"9E",x"A1", -- 0x2308
		x"27",x"C5",x"55",x"96",x"33",x"87",x"9E",x"B5", -- 0x2310
		x"0A",x"6A",x"F0",x"86",x"48",x"8B",x"7C",x"B6", -- 0x2318
		x"83",x"4A",x"54",x"05",x"CA",x"B1",x"87",x"8B", -- 0x2320
		x"2A",x"5C",x"55",x"9F",x"1E",x"74",x"41",x"C4", -- 0x2328
		x"B9",x"16",x"5C",x"EC",x"1D",x"7A",x"A3",x"27", -- 0x2330
		x"64",x"14",x"2D",x"AD",x"1F",x"29",x"E3",x"A2", -- 0x2338
		x"F3",x"B7",x"27",x"BE",x"69",x"AF",x"4A",x"94", -- 0x2340
		x"8B",x"1F",x"B3",x"29",x"13",x"74",x"ED",x"CC", -- 0x2348
		x"8A",x"C9",x"3A",x"27",x"45",x"5D",x"CD",x"A9", -- 0x2350
		x"71",x"FA",x"D6",x"10",x"24",x"3B",x"B2",x"18", -- 0x2358
		x"F2",x"59",x"56",x"DC",x"09",x"20",x"71",x"94", -- 0x2360
		x"BF",x"25",x"BD",x"D2",x"99",x"2C",x"20",x"A3", -- 0x2368
		x"F5",x"5A",x"4A",x"3B",x"B7",x"18",x"65",x"A8", -- 0x2370
		x"13",x"BB",x"38",x"B6",x"76",x"EA",x"4F",x"E9", -- 0x2378
		x"C3",x"A5",x"C6",x"CD",x"46",x"38",x"E1",x"06", -- 0x2380
		x"DC",x"20",x"D8",x"F5",x"4C",x"78",x"19",x"42", -- 0x2388
		x"D2",x"63",x"FD",x"0A",x"7B",x"E2",x"32",x"0E", -- 0x2390
		x"9E",x"6A",x"44",x"95",x"D4",x"93",x"7F",x"99", -- 0x2398
		x"B9",x"46",x"67",x"00",x"FD",x"C8",x"06",x"DA", -- 0x23A0
		x"E8",x"5E",x"50",x"B4",x"D7",x"69",x"F7",x"2A", -- 0x23A8
		x"CC",x"75",x"B4",x"C7",x"58",x"E6",x"D5",x"76", -- 0x23B0
		x"D1",x"99",x"0C",x"A6",x"2E",x"8B",x"40",x"67", -- 0x23B8
		x"51",x"27",x"67",x"4F",x"70",x"EC",x"A9",x"59", -- 0x23C0
		x"4B",x"F9",x"0F",x"A2",x"E2",x"86",x"CD",x"AF", -- 0x23C8
		x"FB",x"02",x"F6",x"D3",x"E8",x"4C",x"C9",x"BA", -- 0x23D0
		x"E6",x"D6",x"E1",x"15",x"E1",x"A1",x"7C",x"B3", -- 0x23D8
		x"C9",x"63",x"82",x"B9",x"50",x"2D",x"13",x"1B", -- 0x23E0
		x"A6",x"A1",x"BE",x"8A",x"A7",x"0C",x"B9",x"23", -- 0x23E8
		x"0E",x"B1",x"F6",x"76",x"FD",x"41",x"B1",x"E4", -- 0x23F0
		x"18",x"93",x"79",x"79",x"35",x"75",x"2D",x"7E", -- 0x23F8
		x"D8",x"B0",x"38",x"A8",x"5D",x"CB",x"C4",x"83", -- 0x2400
		x"EC",x"03",x"0E",x"95",x"0F",x"C8",x"38",x"9C", -- 0x2408
		x"F9",x"AF",x"92",x"F7",x"F0",x"44",x"5D",x"88", -- 0x2410
		x"D7",x"56",x"02",x"8D",x"CC",x"AF",x"8B",x"25", -- 0x2418
		x"60",x"C4",x"CE",x"3D",x"10",x"13",x"C0",x"7C", -- 0x2420
		x"16",x"4F",x"91",x"25",x"97",x"CA",x"41",x"91", -- 0x2428
		x"7A",x"D3",x"09",x"6B",x"19",x"E5",x"F3",x"70", -- 0x2430
		x"3D",x"75",x"7D",x"89",x"25",x"0A",x"AE",x"05", -- 0x2438
		x"4E",x"FC",x"42",x"DD",x"10",x"83",x"5A",x"26", -- 0x2440
		x"D2",x"EC",x"CA",x"6A",x"B7",x"0C",x"7B",x"B1", -- 0x2448
		x"60",x"04",x"1D",x"F8",x"EA",x"90",x"E8",x"A7", -- 0x2450
		x"06",x"67",x"31",x"2C",x"F0",x"5F",x"31",x"3F", -- 0x2458
		x"5D",x"F3",x"9C",x"6D",x"77",x"F6",x"14",x"C9", -- 0x2460
		x"63",x"DE",x"B3",x"1B",x"6B",x"2F",x"CC",x"CB", -- 0x2468
		x"33",x"69",x"C4",x"9D",x"F9",x"AD",x"45",x"80", -- 0x2470
		x"94",x"76",x"AC",x"85",x"D6",x"5D",x"44",x"B3", -- 0x2478
		x"D0",x"E0",x"A0",x"C7",x"58",x"B4",x"91",x"BB", -- 0x2480
		x"14",x"C4",x"57",x"7F",x"73",x"24",x"4B",x"A7", -- 0x2488
		x"0E",x"8F",x"C4",x"08",x"BC",x"0B",x"88",x"D1", -- 0x2490
		x"01",x"B4",x"D6",x"57",x"92",x"1C",x"0B",x"63", -- 0x2498
		x"7C",x"AC",x"AB",x"D4",x"E0",x"3D",x"11",x"F4", -- 0x24A0
		x"82",x"68",x"74",x"F5",x"0C",x"3F",x"1D",x"1A", -- 0x24A8
		x"4E",x"E2",x"A2",x"0C",x"ED",x"AA",x"5D",x"6E", -- 0x24B0
		x"60",x"34",x"C6",x"72",x"50",x"D1",x"55",x"4D", -- 0x24B8
		x"FD",x"01",x"A1",x"DF",x"BE",x"B2",x"D4",x"41", -- 0x24C0
		x"1B",x"4A",x"37",x"28",x"09",x"D4",x"42",x"58", -- 0x24C8
		x"B7",x"E4",x"E3",x"25",x"10",x"41",x"93",x"70", -- 0x24D0
		x"75",x"5A",x"62",x"46",x"AC",x"B7",x"13",x"AA", -- 0x24D8
		x"B9",x"B4",x"8A",x"78",x"68",x"DF",x"B9",x"03", -- 0x24E0
		x"2A",x"70",x"AA",x"B2",x"45",x"6D",x"0B",x"FC", -- 0x24E8
		x"D1",x"6E",x"A1",x"E1",x"2F",x"B5",x"52",x"25", -- 0x24F0
		x"10",x"B4",x"6B",x"3C",x"6D",x"FD",x"E7",x"A6", -- 0x24F8
		x"B2",x"F1",x"1F",x"9A",x"D1",x"D8",x"1E",x"7B", -- 0x2500
		x"C8",x"C8",x"2F",x"0F",x"36",x"B9",x"8B",x"09", -- 0x2508
		x"29",x"AD",x"EA",x"D7",x"63",x"BD",x"FC",x"F2", -- 0x2510
		x"F1",x"68",x"30",x"DE",x"E5",x"18",x"85",x"99", -- 0x2518
		x"89",x"A4",x"B3",x"5C",x"FC",x"D1",x"D7",x"C6", -- 0x2520
		x"1B",x"86",x"55",x"51",x"C0",x"E0",x"D9",x"69", -- 0x2528
		x"8E",x"C5",x"41",x"F1",x"03",x"3F",x"E5",x"F4", -- 0x2530
		x"27",x"95",x"D4",x"0E",x"2D",x"D9",x"27",x"B6", -- 0x2538
		x"7F",x"DA",x"92",x"FB",x"2D",x"EA",x"C2",x"48", -- 0x2540
		x"71",x"18",x"19",x"32",x"79",x"F3",x"9B",x"87", -- 0x2548
		x"39",x"DD",x"7A",x"3C",x"9C",x"DF",x"31",x"C3", -- 0x2550
		x"F4",x"85",x"D1",x"22",x"60",x"F8",x"D8",x"5F", -- 0x2558
		x"54",x"EB",x"5B",x"81",x"D6",x"9E",x"49",x"48", -- 0x2560
		x"B6",x"62",x"FA",x"AF",x"D5",x"16",x"38",x"0F", -- 0x2568
		x"73",x"32",x"CA",x"10",x"91",x"7C",x"D4",x"86", -- 0x2570
		x"02",x"26",x"A8",x"E1",x"20",x"01",x"C0",x"F3", -- 0x2578
		x"EC",x"1D",x"75",x"C3",x"BB",x"3E",x"8C",x"F1", -- 0x2580
		x"20",x"07",x"A2",x"F6",x"1D",x"5A",x"85",x"11", -- 0x2588
		x"8C",x"51",x"21",x"1E",x"CD",x"75",x"24",x"4F", -- 0x2590
		x"9C",x"4C",x"B1",x"3C",x"4D",x"72",x"30",x"BA", -- 0x2598
		x"0F",x"25",x"FD",x"CA",x"E2",x"0A",x"3D",x"03", -- 0x25A0
		x"11",x"DF",x"79",x"AE",x"3A",x"00",x"BF",x"46", -- 0x25A8
		x"D0",x"60",x"E3",x"1E",x"56",x"08",x"EC",x"F2", -- 0x25B0
		x"54",x"9E",x"AE",x"21",x"91",x"5E",x"5B",x"A0", -- 0x25B8
		x"83",x"D9",x"EB",x"66",x"E3",x"29",x"E8",x"75", -- 0x25C0
		x"88",x"63",x"A3",x"C2",x"E2",x"63",x"88",x"33", -- 0x25C8
		x"43",x"6C",x"D0",x"99",x"74",x"BD",x"0C",x"48", -- 0x25D0
		x"DC",x"BA",x"E8",x"6E",x"98",x"C4",x"8E",x"1C", -- 0x25D8
		x"9E",x"7A",x"02",x"02",x"A3",x"6B",x"77",x"2C", -- 0x25E0
		x"4E",x"1B",x"6E",x"B0",x"FD",x"F6",x"E3",x"C1", -- 0x25E8
		x"E2",x"34",x"DA",x"D6",x"F1",x"E7",x"9E",x"4E", -- 0x25F0
		x"22",x"88",x"3C",x"BB",x"4D",x"CB",x"57",x"EB", -- 0x25F8
		x"C5",x"5A",x"6D",x"E9",x"45",x"E5",x"95",x"93", -- 0x2600
		x"80",x"05",x"44",x"FE",x"7B",x"A7",x"C0",x"DE", -- 0x2608
		x"DB",x"9B",x"B5",x"4D",x"03",x"55",x"1C",x"26", -- 0x2610
		x"DD",x"58",x"61",x"AA",x"A3",x"B8",x"16",x"6A", -- 0x2618
		x"92",x"83",x"54",x"D7",x"E8",x"E9",x"6B",x"6A", -- 0x2620
		x"6E",x"2F",x"E8",x"6A",x"56",x"29",x"49",x"B1", -- 0x2628
		x"44",x"FE",x"7F",x"48",x"D3",x"9B",x"ED",x"31", -- 0x2630
		x"F3",x"4F",x"DB",x"98",x"08",x"71",x"82",x"9B", -- 0x2638
		x"F5",x"D6",x"F2",x"DE",x"40",x"DE",x"C8",x"AF", -- 0x2640
		x"0E",x"31",x"1A",x"E4",x"5A",x"E2",x"96",x"9F", -- 0x2648
		x"E1",x"16",x"E7",x"B6",x"B1",x"D5",x"67",x"26", -- 0x2650
		x"A4",x"44",x"3E",x"AC",x"B5",x"C0",x"C7",x"2B", -- 0x2658
		x"17",x"BB",x"8A",x"57",x"9A",x"D2",x"86",x"28", -- 0x2660
		x"05",x"20",x"0D",x"5F",x"03",x"24",x"FE",x"65", -- 0x2668
		x"B9",x"66",x"9B",x"EB",x"BB",x"03",x"12",x"60", -- 0x2670
		x"C6",x"50",x"8D",x"FC",x"90",x"D4",x"28",x"A7", -- 0x2678
		x"90",x"32",x"FE",x"AA",x"06",x"86",x"53",x"0B", -- 0x2680
		x"A6",x"DF",x"6A",x"2A",x"83",x"E9",x"8F",x"3E", -- 0x2688
		x"CF",x"2B",x"2A",x"8C",x"2E",x"BB",x"6C",x"F5", -- 0x2690
		x"0C",x"F9",x"F2",x"1C",x"4F",x"9A",x"C3",x"DF", -- 0x2698
		x"CD",x"C2",x"0B",x"D3",x"C8",x"5E",x"5E",x"EF", -- 0x26A0
		x"BD",x"C8",x"1A",x"42",x"32",x"A9",x"80",x"03", -- 0x26A8
		x"D4",x"2A",x"0F",x"82",x"E5",x"7B",x"F7",x"71", -- 0x26B0
		x"F5",x"EA",x"8D",x"45",x"06",x"51",x"A4",x"D3", -- 0x26B8
		x"93",x"AF",x"27",x"5D",x"8D",x"85",x"4D",x"CB", -- 0x26C0
		x"4E",x"E6",x"0E",x"01",x"90",x"0E",x"04",x"E4", -- 0x26C8
		x"38",x"13",x"E6",x"1E",x"0E",x"DF",x"0F",x"04", -- 0x26D0
		x"4A",x"9C",x"C8",x"50",x"ED",x"6E",x"A3",x"81", -- 0x26D8
		x"9D",x"CA",x"5E",x"AB",x"50",x"2B",x"77",x"1F", -- 0x26E0
		x"12",x"05",x"20",x"22",x"92",x"A3",x"07",x"CA", -- 0x26E8
		x"36",x"6E",x"68",x"C3",x"4E",x"77",x"C8",x"98", -- 0x26F0
		x"93",x"11",x"69",x"01",x"7F",x"0D",x"02",x"9D", -- 0x26F8
		x"D8",x"61",x"C8",x"29",x"8C",x"BF",x"C7",x"1F", -- 0x2700
		x"C4",x"67",x"41",x"57",x"0B",x"C8",x"A1",x"C0", -- 0x2708
		x"37",x"89",x"85",x"85",x"80",x"CD",x"9D",x"14", -- 0x2710
		x"DE",x"86",x"15",x"DE",x"94",x"17",x"7C",x"EC", -- 0x2718
		x"F7",x"45",x"95",x"85",x"05",x"5E",x"A4",x"49", -- 0x2720
		x"C5",x"65",x"20",x"51",x"2E",x"41",x"12",x"65", -- 0x2728
		x"CA",x"97",x"6A",x"4B",x"65",x"09",x"DE",x"45", -- 0x2730
		x"0F",x"F3",x"24",x"A3",x"8A",x"20",x"90",x"83", -- 0x2738
		x"65",x"27",x"88",x"E9",x"05",x"AC",x"B2",x"CA", -- 0x2740
		x"12",x"D2",x"1C",x"41",x"14",x"2F",x"A6",x"5E", -- 0x2748
		x"46",x"12",x"29",x"AC",x"9A",x"08",x"71",x"A9", -- 0x2750
		x"7B",x"15",x"CD",x"85",x"35",x"DD",x"09",x"1A", -- 0x2758
		x"05",x"91",x"83",x"89",x"3E",x"36",x"55",x"D0", -- 0x2760
		x"88",x"F0",x"12",x"1C",x"9F",x"38",x"7A",x"E6", -- 0x2768
		x"C9",x"23",x"13",x"64",x"2B",x"84",x"8E",x"26", -- 0x2770
		x"99",x"DB",x"AB",x"4E",x"B9",x"35",x"E7",x"3F", -- 0x2778
		x"C6",x"6B",x"C8",x"85",x"21",x"9D",x"56",x"A9", -- 0x2780
		x"8F",x"E7",x"C5",x"2F",x"20",x"BF",x"16",x"EA", -- 0x2788
		x"E2",x"29",x"CE",x"8D",x"2D",x"DC",x"33",x"46", -- 0x2790
		x"B8",x"DE",x"94",x"73",x"14",x"FB",x"32",x"5B", -- 0x2798
		x"67",x"FA",x"60",x"88",x"99",x"36",x"B1",x"A8", -- 0x27A0
		x"9D",x"77",x"D7",x"BD",x"B6",x"6E",x"28",x"99", -- 0x27A8
		x"17",x"F7",x"A6",x"45",x"54",x"D9",x"0B",x"0E", -- 0x27B0
		x"B9",x"A0",x"01",x"4D",x"1C",x"B2",x"28",x"84", -- 0x27B8
		x"AD",x"08",x"8C",x"C6",x"3E",x"3F",x"6F",x"DB", -- 0x27C0
		x"36",x"C7",x"1A",x"ED",x"36",x"42",x"07",x"CC", -- 0x27C8
		x"B9",x"AE",x"12",x"0F",x"88",x"1E",x"9C",x"C1", -- 0x27D0
		x"3E",x"1D",x"8F",x"D9",x"CF",x"B7",x"5E",x"FC", -- 0x27D8
		x"40",x"6B",x"C4",x"FD",x"2A",x"B3",x"5A",x"DF", -- 0x27E0
		x"FA",x"74",x"CD",x"B0",x"36",x"55",x"7E",x"70", -- 0x27E8
		x"04",x"10",x"7F",x"0C",x"AD",x"9B",x"CE",x"6B", -- 0x27F0
		x"B8",x"DD",x"46",x"08",x"15",x"24",x"05",x"55", -- 0x27F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2808
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2810
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2820
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2828
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2830
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2840
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2850
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2858
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2860
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2868
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2870
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2878
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2880
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2888
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2890
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2898
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x28F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2900
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2908
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2910
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2918
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2920
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2928
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2930
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2938
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2940
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2948
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2950
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2958
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2960
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2968
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2970
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2978
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2980
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2988
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2990
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2998
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x29F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2A98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2AF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x2FF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3000
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3008
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3010
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3018
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3020
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3028
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3030
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3038
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3040
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3048
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3050
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3058
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3060
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3068
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3070
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3078
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3080
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3088
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3090
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3098
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x30F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3100
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3108
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3110
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3118
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3120
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3128
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3130
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3138
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3140
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3148
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3150
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3158
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3160
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3168
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3170
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3178
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3180
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3188
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3190
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3198
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x31F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3200
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3208
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3210
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3218
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3220
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3228
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3230
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3238
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3240
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3248
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3250
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3258
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3260
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3268
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3270
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3278
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3280
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3288
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3290
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3298
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x32F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3300
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3308
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3310
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3318
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3320
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3328
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3330
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3338
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3340
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3348
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3350
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3358
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3360
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3368
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3370
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3378
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3380
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3388
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3390
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3398
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x33F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3400
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3408
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3410
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3418
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3420
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3430
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3438
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3440
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3448
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3450
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3458
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3460
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3468
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3470
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3478
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3480
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3488
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3490
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3498
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x34F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3500
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3508
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3510
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3518
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3520
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3528
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3530
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3538
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3540
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3548
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3550
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3558
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3560
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3568
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3570
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3578
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3580
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3588
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3590
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3598
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x35F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3600
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3608
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3610
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3618
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3620
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3628
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3630
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3638
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3640
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3648
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3650
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3658
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3660
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3668
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3670
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3678
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3680
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3688
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3690
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3698
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x36F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3700
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3708
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3710
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3718
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3720
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3728
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3730
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3738
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3740
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3748
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3750
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3758
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3760
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3768
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3770
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3778
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3780
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3788
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3790
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3798
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x37F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3800
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3808
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3810
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3818
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3820
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3828
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3830
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3838
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3840
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3848
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3850
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3858
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3860
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3868
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3870
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3878
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3880
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3888
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3890
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3898
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x38F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3900
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3908
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3910
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3918
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3920
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3928
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3930
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3938
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3940
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3948
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3950
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3958
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3960
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3968
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3970
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3978
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3980
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3988
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3990
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3998
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39A8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x39F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3A98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3AF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3B98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3BF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3C98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3CF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3D98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3DF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3E98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3ED0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3ED8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3EF8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F00
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F08
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F10
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F18
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F20
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F28
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F30
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F38
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F40
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F48
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F50
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F58
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F60
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F68
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F70
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F78
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F80
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F88
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F90
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3F98
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FA8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FB8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FC8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FD8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FE8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x3FF0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x3FF8
	);
	attribute ram_style : string;
	attribute ram_style of ROM : signal is "block";

begin

	p_rom : process(CLK,ADDR)
	begin
		if (rising_edge(CLK)) then
			DATA <= ROM(to_integer(unsigned(ADDR)));
		 end if;
	end process;
end RTL;
