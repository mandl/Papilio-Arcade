-- generated with romgen v3.04 by MikeJ
-- dummy rom. random rom data. avoid map to optimise this rom away;
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

--library UNISIM;
	--use UNISIM.Vcomponents.all;

entity INVADERS_ROM is
port (
	CLK  : in  std_logic;
	ADDR : in  std_logic_vector(12 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of INVADERS_ROM is


	type ROM_ARRAY is array(0 to 8191) of std_logic_vector(7 downto 0);
	signal ROM : ROM_ARRAY := (
		x"FB",x"DE",x"3B",x"A4",x"C4",x"F1",x"65",x"6E", -- 0x0000
		x"97",x"81",x"E9",x"8A",x"A4",x"17",x"5B",x"A2", -- 0x0008
		x"20",x"B8",x"63",x"F2",x"44",x"2D",x"4F",x"42", -- 0x0010
		x"79",x"9B",x"A3",x"A5",x"4B",x"0B",x"09",x"47", -- 0x0018
		x"E9",x"C3",x"6C",x"AF",x"35",x"D1",x"9D",x"CD", -- 0x0020
		x"D3",x"88",x"D7",x"F7",x"1F",x"33",x"9A",x"40", -- 0x0028
		x"6B",x"7E",x"B2",x"B0",x"AB",x"03",x"F2",x"A4", -- 0x0030
		x"1E",x"17",x"4A",x"69",x"22",x"D2",x"30",x"8C", -- 0x0038
		x"96",x"9C",x"3C",x"CC",x"EE",x"D9",x"1A",x"42", -- 0x0040
		x"E1",x"F1",x"3A",x"81",x"25",x"55",x"C1",x"91", -- 0x0048
		x"D3",x"74",x"C1",x"FE",x"F6",x"B4",x"23",x"15", -- 0x0050
		x"4B",x"EC",x"7E",x"6E",x"C0",x"2F",x"FA",x"D6", -- 0x0058
		x"4B",x"B6",x"23",x"3A",x"10",x"3D",x"7C",x"F2", -- 0x0060
		x"AE",x"37",x"74",x"54",x"8C",x"B5",x"65",x"DF", -- 0x0068
		x"A9",x"27",x"5E",x"A1",x"5B",x"81",x"B6",x"A7", -- 0x0070
		x"ED",x"B5",x"16",x"AE",x"64",x"11",x"06",x"AF", -- 0x0078
		x"47",x"A8",x"EA",x"57",x"E6",x"E6",x"C9",x"15", -- 0x0080
		x"9D",x"BD",x"69",x"2A",x"73",x"CE",x"89",x"9D", -- 0x0088
		x"F5",x"E7",x"3F",x"52",x"E8",x"75",x"F9",x"D7", -- 0x0090
		x"AA",x"8F",x"86",x"0F",x"20",x"0C",x"3F",x"67", -- 0x0098
		x"B5",x"A9",x"BE",x"1C",x"90",x"09",x"B0",x"AE", -- 0x00A0
		x"C6",x"1B",x"D8",x"3B",x"69",x"E2",x"58",x"60", -- 0x00A8
		x"CA",x"97",x"32",x"B4",x"8C",x"AB",x"8C",x"38", -- 0x00B0
		x"3B",x"92",x"C6",x"DA",x"1F",x"06",x"42",x"D4", -- 0x00B8
		x"AF",x"80",x"70",x"C0",x"89",x"21",x"6F",x"51", -- 0x00C0
		x"BB",x"C7",x"0C",x"26",x"2A",x"64",x"86",x"F5", -- 0x00C8
		x"7B",x"38",x"2A",x"08",x"E3",x"B6",x"BF",x"9E", -- 0x00D0
		x"C8",x"07",x"79",x"E7",x"0D",x"3B",x"3C",x"3D", -- 0x00D8
		x"BB",x"2C",x"7D",x"C5",x"CD",x"6C",x"17",x"89", -- 0x00E0
		x"34",x"A2",x"AF",x"5F",x"86",x"B5",x"D4",x"02", -- 0x00E8
		x"ED",x"FE",x"89",x"51",x"35",x"4A",x"6F",x"7D", -- 0x00F0
		x"51",x"E8",x"E5",x"DD",x"24",x"A1",x"9A",x"60", -- 0x00F8
		x"4E",x"18",x"26",x"1C",x"84",x"BC",x"A5",x"39", -- 0x0100
		x"5F",x"D5",x"18",x"E5",x"0B",x"EC",x"67",x"79", -- 0x0108
		x"6B",x"F0",x"CA",x"20",x"BA",x"BA",x"1D",x"8B", -- 0x0110
		x"A3",x"03",x"E9",x"48",x"25",x"84",x"28",x"73", -- 0x0118
		x"9D",x"4E",x"8F",x"A1",x"8A",x"B4",x"DA",x"E9", -- 0x0120
		x"8A",x"F2",x"4F",x"16",x"5F",x"B6",x"8F",x"4A", -- 0x0128
		x"27",x"D9",x"6A",x"E2",x"94",x"88",x"ED",x"B8", -- 0x0130
		x"0B",x"D7",x"80",x"30",x"DC",x"A8",x"A3",x"7A", -- 0x0138
		x"76",x"B2",x"1C",x"01",x"68",x"77",x"6A",x"72", -- 0x0140
		x"6A",x"B9",x"88",x"4A",x"EF",x"97",x"94",x"17", -- 0x0148
		x"72",x"7F",x"79",x"07",x"87",x"68",x"3F",x"92", -- 0x0150
		x"BF",x"BF",x"43",x"9C",x"E7",x"66",x"96",x"5E", -- 0x0158
		x"99",x"33",x"5F",x"02",x"AA",x"C9",x"F3",x"15", -- 0x0160
		x"03",x"FC",x"DE",x"F2",x"14",x"74",x"8A",x"86", -- 0x0168
		x"F3",x"04",x"0E",x"FA",x"EB",x"4D",x"0D",x"AC", -- 0x0170
		x"8D",x"50",x"C8",x"75",x"37",x"60",x"D4",x"D0", -- 0x0178
		x"93",x"B3",x"52",x"3E",x"FD",x"C5",x"D2",x"01", -- 0x0180
		x"C2",x"B2",x"74",x"D7",x"A6",x"FE",x"DD",x"1A", -- 0x0188
		x"03",x"6B",x"15",x"EF",x"B9",x"22",x"1C",x"47", -- 0x0190
		x"F2",x"E4",x"3C",x"2A",x"45",x"11",x"FA",x"58", -- 0x0198
		x"45",x"CC",x"96",x"43",x"92",x"E9",x"44",x"D5", -- 0x01A0
		x"9C",x"B8",x"2D",x"43",x"37",x"0B",x"DC",x"3B", -- 0x01A8
		x"77",x"F1",x"AA",x"B0",x"14",x"46",x"77",x"07", -- 0x01B0
		x"AA",x"B3",x"B0",x"70",x"45",x"2B",x"C8",x"8A", -- 0x01B8
		x"F7",x"60",x"CD",x"8B",x"C9",x"91",x"61",x"66", -- 0x01C0
		x"CA",x"8E",x"29",x"02",x"19",x"06",x"BC",x"90", -- 0x01C8
		x"77",x"67",x"C0",x"8B",x"2D",x"38",x"13",x"D8", -- 0x01D0
		x"6C",x"C3",x"49",x"B1",x"EF",x"12",x"3C",x"E7", -- 0x01D8
		x"F1",x"89",x"F2",x"BB",x"9A",x"D3",x"A1",x"65", -- 0x01E0
		x"E1",x"4A",x"E7",x"FB",x"50",x"A4",x"0C",x"47", -- 0x01E8
		x"8C",x"CD",x"D3",x"B9",x"85",x"66",x"92",x"F1", -- 0x01F0
		x"A9",x"DB",x"A3",x"99",x"6E",x"5F",x"02",x"60", -- 0x01F8
		x"68",x"74",x"9C",x"04",x"49",x"3E",x"E8",x"2B", -- 0x0200
		x"89",x"D0",x"A6",x"59",x"F5",x"B3",x"A1",x"82", -- 0x0208
		x"01",x"F4",x"BB",x"86",x"5B",x"CE",x"F8",x"84", -- 0x0210
		x"AA",x"1C",x"9E",x"98",x"7C",x"A0",x"F9",x"64", -- 0x0218
		x"94",x"16",x"68",x"DD",x"54",x"D1",x"89",x"5D", -- 0x0220
		x"22",x"30",x"B7",x"18",x"63",x"D8",x"1A",x"64", -- 0x0228
		x"CD",x"D6",x"6B",x"A8",x"A5",x"64",x"2D",x"CF", -- 0x0230
		x"80",x"CB",x"E8",x"7C",x"EB",x"E2",x"E1",x"01", -- 0x0238
		x"F8",x"C9",x"5E",x"CC",x"9B",x"E7",x"2B",x"BE", -- 0x0240
		x"98",x"62",x"56",x"7B",x"3B",x"71",x"60",x"88", -- 0x0248
		x"C7",x"CB",x"31",x"EC",x"AF",x"DD",x"3C",x"30", -- 0x0250
		x"2A",x"25",x"2D",x"95",x"87",x"8E",x"96",x"00", -- 0x0258
		x"D7",x"75",x"CD",x"74",x"5D",x"78",x"B2",x"75", -- 0x0260
		x"DA",x"88",x"F1",x"16",x"79",x"D1",x"9E",x"41", -- 0x0268
		x"9D",x"4F",x"AD",x"4D",x"AC",x"EA",x"FC",x"56", -- 0x0270
		x"8F",x"2A",x"6C",x"18",x"38",x"82",x"97",x"11", -- 0x0278
		x"F7",x"65",x"05",x"D5",x"5D",x"37",x"4B",x"38", -- 0x0280
		x"BF",x"BC",x"CD",x"3A",x"8E",x"EB",x"FA",x"AB", -- 0x0288
		x"3B",x"29",x"78",x"68",x"93",x"76",x"3E",x"23", -- 0x0290
		x"20",x"AA",x"BA",x"59",x"AD",x"53",x"E9",x"A5", -- 0x0298
		x"38",x"EE",x"7B",x"96",x"26",x"47",x"4E",x"65", -- 0x02A0
		x"83",x"1D",x"9F",x"92",x"09",x"1B",x"BD",x"C4", -- 0x02A8
		x"44",x"37",x"AC",x"D7",x"AD",x"6A",x"7A",x"4D", -- 0x02B0
		x"95",x"36",x"26",x"43",x"09",x"10",x"E8",x"C0", -- 0x02B8
		x"FE",x"E4",x"57",x"A4",x"AB",x"26",x"0B",x"AE", -- 0x02C0
		x"C2",x"2A",x"C0",x"CB",x"45",x"7F",x"10",x"09", -- 0x02C8
		x"B6",x"3C",x"60",x"E3",x"A7",x"DB",x"B0",x"3D", -- 0x02D0
		x"91",x"D7",x"80",x"1A",x"E7",x"E8",x"DA",x"67", -- 0x02D8
		x"4D",x"B2",x"0C",x"F8",x"D8",x"96",x"28",x"9B", -- 0x02E0
		x"C1",x"E8",x"E6",x"86",x"68",x"77",x"10",x"9E", -- 0x02E8
		x"B3",x"70",x"02",x"DA",x"CB",x"B3",x"97",x"5D", -- 0x02F0
		x"8B",x"18",x"77",x"F2",x"81",x"53",x"5A",x"CE", -- 0x02F8
		x"06",x"E6",x"48",x"5E",x"FC",x"70",x"79",x"BE", -- 0x0300
		x"D8",x"60",x"C5",x"42",x"57",x"D5",x"60",x"8B", -- 0x0308
		x"46",x"63",x"66",x"13",x"17",x"FE",x"EF",x"22", -- 0x0310
		x"96",x"E7",x"15",x"18",x"BA",x"EF",x"67",x"40", -- 0x0318
		x"56",x"2F",x"9E",x"53",x"1F",x"18",x"92",x"F7", -- 0x0320
		x"F7",x"58",x"B9",x"CF",x"AD",x"1B",x"5B",x"F3", -- 0x0328
		x"FD",x"C1",x"86",x"94",x"40",x"F6",x"B6",x"D7", -- 0x0330
		x"DE",x"4B",x"6F",x"19",x"BA",x"56",x"59",x"11", -- 0x0338
		x"05",x"F7",x"E4",x"24",x"8F",x"77",x"1D",x"07", -- 0x0340
		x"4F",x"56",x"D6",x"FC",x"F0",x"32",x"70",x"EE", -- 0x0348
		x"74",x"F7",x"83",x"34",x"6E",x"B9",x"0C",x"CC", -- 0x0350
		x"06",x"FB",x"E5",x"C0",x"D1",x"3F",x"52",x"D7", -- 0x0358
		x"B6",x"37",x"FB",x"C5",x"AE",x"98",x"CC",x"FD", -- 0x0360
		x"6F",x"24",x"FA",x"60",x"D5",x"6B",x"50",x"4A", -- 0x0368
		x"E2",x"53",x"FE",x"D0",x"0E",x"8A",x"9D",x"14", -- 0x0370
		x"86",x"83",x"54",x"D8",x"42",x"A6",x"B0",x"F8", -- 0x0378
		x"DD",x"2C",x"BE",x"8C",x"45",x"0C",x"0A",x"B4", -- 0x0380
		x"AF",x"05",x"15",x"85",x"F0",x"E4",x"50",x"53", -- 0x0388
		x"39",x"4F",x"25",x"47",x"D9",x"C2",x"DA",x"E0", -- 0x0390
		x"C6",x"2F",x"B9",x"09",x"D6",x"E9",x"03",x"B4", -- 0x0398
		x"16",x"41",x"C1",x"DA",x"4D",x"CB",x"0F",x"7C", -- 0x03A0
		x"51",x"A4",x"03",x"42",x"89",x"53",x"95",x"42", -- 0x03A8
		x"22",x"3A",x"09",x"FB",x"FD",x"E3",x"5C",x"C4", -- 0x03B0
		x"93",x"16",x"4D",x"6A",x"00",x"50",x"9E",x"96", -- 0x03B8
		x"12",x"DF",x"F0",x"5F",x"2C",x"01",x"DC",x"7D", -- 0x03C0
		x"A5",x"5F",x"3F",x"AE",x"32",x"54",x"F1",x"54", -- 0x03C8
		x"8F",x"7A",x"CF",x"0D",x"5F",x"2D",x"D1",x"F2", -- 0x03D0
		x"C2",x"9E",x"DC",x"43",x"EF",x"FA",x"59",x"02", -- 0x03D8
		x"5B",x"4A",x"E0",x"87",x"CA",x"3D",x"84",x"70", -- 0x03E0
		x"9C",x"C3",x"9F",x"4E",x"18",x"11",x"A2",x"27", -- 0x03E8
		x"8B",x"F2",x"34",x"EA",x"9F",x"85",x"5D",x"62", -- 0x03F0
		x"25",x"B9",x"A5",x"15",x"35",x"FE",x"96",x"90", -- 0x03F8
		x"4A",x"F6",x"97",x"15",x"35",x"1C",x"06",x"51", -- 0x0400
		x"5F",x"25",x"20",x"77",x"36",x"C2",x"9F",x"C1", -- 0x0408
		x"35",x"D3",x"2D",x"D4",x"D9",x"0A",x"38",x"FE", -- 0x0410
		x"C4",x"5D",x"93",x"79",x"5D",x"2A",x"89",x"27", -- 0x0418
		x"21",x"21",x"BB",x"D5",x"BC",x"41",x"A7",x"1C", -- 0x0420
		x"66",x"C7",x"93",x"1C",x"0A",x"B2",x"DE",x"40", -- 0x0428
		x"07",x"8B",x"94",x"E0",x"95",x"CC",x"DF",x"D9", -- 0x0430
		x"AA",x"73",x"53",x"87",x"1D",x"DC",x"2E",x"BD", -- 0x0438
		x"7D",x"E9",x"94",x"3A",x"AB",x"3C",x"56",x"91", -- 0x0440
		x"83",x"6A",x"AE",x"8D",x"1D",x"0D",x"4D",x"A3", -- 0x0448
		x"98",x"E2",x"04",x"2E",x"2F",x"E3",x"88",x"D9", -- 0x0450
		x"D6",x"DB",x"61",x"73",x"39",x"8F",x"32",x"36", -- 0x0458
		x"F9",x"46",x"71",x"25",x"02",x"C7",x"B6",x"85", -- 0x0460
		x"B1",x"E4",x"92",x"CF",x"F1",x"E0",x"F2",x"0A", -- 0x0468
		x"C3",x"F7",x"B8",x"72",x"5B",x"41",x"4D",x"B2", -- 0x0470
		x"9C",x"2E",x"26",x"55",x"3E",x"58",x"8C",x"38", -- 0x0478
		x"9E",x"FD",x"DC",x"A0",x"45",x"13",x"A5",x"F7", -- 0x0480
		x"F8",x"39",x"47",x"6A",x"1A",x"3A",x"75",x"5D", -- 0x0488
		x"B1",x"AD",x"CF",x"0E",x"EE",x"9C",x"C0",x"0B", -- 0x0490
		x"CB",x"66",x"61",x"0A",x"BF",x"6D",x"C1",x"DD", -- 0x0498
		x"6B",x"1E",x"FE",x"30",x"31",x"24",x"A7",x"A9", -- 0x04A0
		x"5D",x"6E",x"15",x"F6",x"29",x"0A",x"54",x"DA", -- 0x04A8
		x"B7",x"A4",x"68",x"26",x"41",x"29",x"B0",x"8C", -- 0x04B0
		x"90",x"12",x"16",x"CF",x"7F",x"57",x"2D",x"6A", -- 0x04B8
		x"75",x"AB",x"1B",x"27",x"D0",x"C2",x"D0",x"2E", -- 0x04C0
		x"32",x"65",x"A5",x"5B",x"EE",x"F9",x"B5",x"26", -- 0x04C8
		x"1E",x"1F",x"CB",x"DF",x"C7",x"7D",x"6C",x"D7", -- 0x04D0
		x"0F",x"03",x"A7",x"0F",x"5A",x"55",x"F8",x"50", -- 0x04D8
		x"01",x"14",x"F6",x"D1",x"57",x"C7",x"80",x"09", -- 0x04E0
		x"AD",x"26",x"E3",x"1C",x"9F",x"99",x"C2",x"3E", -- 0x04E8
		x"B8",x"8E",x"1E",x"01",x"8B",x"0A",x"D8",x"9B", -- 0x04F0
		x"0D",x"01",x"2A",x"E7",x"56",x"23",x"38",x"57", -- 0x04F8
		x"38",x"2F",x"A9",x"8F",x"76",x"A9",x"18",x"A3", -- 0x0500
		x"4F",x"FB",x"40",x"6E",x"95",x"03",x"AC",x"CE", -- 0x0508
		x"11",x"4A",x"CF",x"1D",x"55",x"A8",x"38",x"62", -- 0x0510
		x"29",x"62",x"4A",x"7F",x"85",x"02",x"57",x"3D", -- 0x0518
		x"B0",x"80",x"CC",x"28",x"A9",x"E4",x"4B",x"F8", -- 0x0520
		x"60",x"8B",x"E6",x"F6",x"0E",x"94",x"45",x"9F", -- 0x0528
		x"5E",x"15",x"BC",x"B3",x"3D",x"F4",x"96",x"67", -- 0x0530
		x"57",x"60",x"66",x"5C",x"63",x"BD",x"9A",x"14", -- 0x0538
		x"BD",x"E6",x"BB",x"67",x"4C",x"87",x"60",x"AC", -- 0x0540
		x"13",x"48",x"23",x"A1",x"5C",x"68",x"41",x"BA", -- 0x0548
		x"FC",x"FD",x"EE",x"BA",x"F2",x"85",x"22",x"C9", -- 0x0550
		x"E5",x"08",x"26",x"C8",x"C6",x"40",x"DD",x"84", -- 0x0558
		x"28",x"19",x"EC",x"74",x"A0",x"CC",x"A0",x"34", -- 0x0560
		x"94",x"C4",x"D5",x"70",x"2D",x"17",x"2C",x"2B", -- 0x0568
		x"94",x"9A",x"E5",x"07",x"20",x"87",x"50",x"85", -- 0x0570
		x"8F",x"F5",x"4F",x"D5",x"37",x"2D",x"DA",x"5F", -- 0x0578
		x"C5",x"47",x"53",x"67",x"93",x"73",x"1B",x"29", -- 0x0580
		x"38",x"F0",x"99",x"E5",x"87",x"45",x"90",x"1C", -- 0x0588
		x"5F",x"76",x"A2",x"7F",x"7D",x"F2",x"85",x"8C", -- 0x0590
		x"E8",x"D4",x"E2",x"20",x"81",x"BD",x"FE",x"47", -- 0x0598
		x"84",x"D1",x"2E",x"18",x"46",x"49",x"C0",x"7E", -- 0x05A0
		x"B9",x"DA",x"64",x"41",x"9F",x"F4",x"DC",x"00", -- 0x05A8
		x"EA",x"FE",x"FE",x"E7",x"F1",x"84",x"F4",x"DB", -- 0x05B0
		x"59",x"D7",x"7B",x"DA",x"15",x"FA",x"A2",x"99", -- 0x05B8
		x"CC",x"D0",x"31",x"13",x"9A",x"F2",x"12",x"54", -- 0x05C0
		x"4D",x"F5",x"16",x"EC",x"6B",x"72",x"EC",x"D5", -- 0x05C8
		x"72",x"6C",x"BE",x"64",x"F0",x"B3",x"BF",x"CA", -- 0x05D0
		x"0B",x"BB",x"A5",x"20",x"B6",x"C7",x"39",x"83", -- 0x05D8
		x"99",x"6A",x"17",x"B3",x"DC",x"29",x"08",x"A9", -- 0x05E0
		x"9E",x"9D",x"97",x"0A",x"11",x"04",x"E0",x"83", -- 0x05E8
		x"70",x"1F",x"67",x"E1",x"D2",x"A7",x"AC",x"5D", -- 0x05F0
		x"63",x"D1",x"7D",x"99",x"9A",x"36",x"9C",x"B3", -- 0x05F8
		x"20",x"B3",x"67",x"7D",x"5C",x"EE",x"27",x"7B", -- 0x0600
		x"8D",x"BE",x"85",x"1E",x"43",x"66",x"A1",x"33", -- 0x0608
		x"85",x"88",x"15",x"D7",x"AF",x"C1",x"35",x"92", -- 0x0610
		x"94",x"32",x"2C",x"AE",x"68",x"C9",x"62",x"09", -- 0x0618
		x"FC",x"C9",x"86",x"D9",x"B8",x"AD",x"55",x"C5", -- 0x0620
		x"EC",x"DA",x"E3",x"30",x"C1",x"05",x"63",x"C6", -- 0x0628
		x"0E",x"F8",x"1F",x"BD",x"BA",x"54",x"51",x"CE", -- 0x0630
		x"07",x"FC",x"FC",x"EE",x"C6",x"5F",x"F7",x"44", -- 0x0638
		x"A8",x"FD",x"9D",x"E1",x"AC",x"F2",x"A7",x"19", -- 0x0640
		x"4D",x"0C",x"C8",x"0F",x"11",x"AB",x"56",x"1F", -- 0x0648
		x"A4",x"75",x"DD",x"DF",x"49",x"AE",x"2E",x"50", -- 0x0650
		x"AB",x"2C",x"40",x"F2",x"8B",x"B7",x"B6",x"B4", -- 0x0658
		x"B6",x"54",x"96",x"E2",x"47",x"BD",x"FB",x"14", -- 0x0660
		x"C9",x"C4",x"A3",x"DB",x"70",x"F9",x"7A",x"95", -- 0x0668
		x"6F",x"D7",x"75",x"B8",x"86",x"A3",x"89",x"B2", -- 0x0670
		x"4F",x"49",x"25",x"5B",x"01",x"DB",x"10",x"37", -- 0x0678
		x"AF",x"A6",x"99",x"F6",x"E3",x"95",x"8A",x"AE", -- 0x0680
		x"D9",x"2E",x"8A",x"CA",x"28",x"84",x"60",x"17", -- 0x0688
		x"5D",x"55",x"50",x"E3",x"78",x"D9",x"16",x"C8", -- 0x0690
		x"23",x"3B",x"24",x"A3",x"96",x"34",x"5B",x"46", -- 0x0698
		x"5A",x"F4",x"BC",x"3E",x"0B",x"48",x"6C",x"E4", -- 0x06A0
		x"76",x"F6",x"2F",x"1F",x"7C",x"0F",x"36",x"59", -- 0x06A8
		x"64",x"86",x"3D",x"DD",x"DF",x"D3",x"26",x"82", -- 0x06B0
		x"0F",x"4A",x"A6",x"A6",x"FD",x"02",x"EC",x"58", -- 0x06B8
		x"F6",x"AA",x"16",x"81",x"F2",x"83",x"E6",x"E8", -- 0x06C0
		x"F9",x"16",x"08",x"F5",x"26",x"BE",x"4F",x"0A", -- 0x06C8
		x"C4",x"0D",x"67",x"A5",x"E0",x"8D",x"28",x"6F", -- 0x06D0
		x"D7",x"CE",x"16",x"55",x"50",x"83",x"AD",x"48", -- 0x06D8
		x"2E",x"44",x"49",x"A0",x"47",x"30",x"09",x"41", -- 0x06E0
		x"47",x"12",x"B7",x"EC",x"50",x"86",x"F6",x"15", -- 0x06E8
		x"93",x"DE",x"BA",x"F3",x"6C",x"63",x"64",x"C4", -- 0x06F0
		x"32",x"7A",x"1A",x"83",x"FD",x"48",x"4B",x"AB", -- 0x06F8
		x"8C",x"94",x"CB",x"53",x"45",x"D5",x"94",x"0C", -- 0x0700
		x"67",x"CB",x"F8",x"37",x"53",x"6F",x"4C",x"66", -- 0x0708
		x"4E",x"08",x"5B",x"3B",x"EA",x"BF",x"00",x"1D", -- 0x0710
		x"B9",x"1A",x"20",x"38",x"62",x"EA",x"63",x"6E", -- 0x0718
		x"00",x"30",x"C1",x"45",x"85",x"D6",x"51",x"6C", -- 0x0720
		x"A2",x"C9",x"A3",x"75",x"B8",x"EF",x"DC",x"08", -- 0x0728
		x"77",x"38",x"C2",x"62",x"77",x"C2",x"00",x"31", -- 0x0730
		x"5C",x"9F",x"E8",x"BF",x"8B",x"4D",x"AD",x"0B", -- 0x0738
		x"7D",x"EF",x"50",x"82",x"C6",x"21",x"EE",x"E8", -- 0x0740
		x"6A",x"12",x"5F",x"23",x"02",x"BB",x"AA",x"F9", -- 0x0748
		x"F3",x"6D",x"DB",x"EA",x"AF",x"DB",x"9B",x"0D", -- 0x0750
		x"FB",x"85",x"4C",x"07",x"D2",x"F9",x"12",x"CF", -- 0x0758
		x"E9",x"E1",x"52",x"30",x"82",x"C0",x"1A",x"EC", -- 0x0760
		x"D2",x"79",x"10",x"D4",x"35",x"3B",x"4E",x"A8", -- 0x0768
		x"A8",x"2B",x"13",x"59",x"86",x"AE",x"66",x"02", -- 0x0770
		x"34",x"32",x"09",x"86",x"AB",x"1B",x"56",x"96", -- 0x0778
		x"FC",x"A8",x"C6",x"FE",x"69",x"60",x"EB",x"BB", -- 0x0780
		x"59",x"7C",x"11",x"0E",x"B7",x"5F",x"36",x"60", -- 0x0788
		x"0A",x"49",x"39",x"11",x"78",x"1F",x"13",x"2C", -- 0x0790
		x"51",x"1D",x"B3",x"FD",x"B7",x"89",x"14",x"B5", -- 0x0798
		x"B2",x"5A",x"34",x"1C",x"BB",x"21",x"58",x"94", -- 0x07A0
		x"9D",x"69",x"A3",x"55",x"C8",x"D9",x"35",x"D3", -- 0x07A8
		x"24",x"EE",x"64",x"9C",x"0E",x"77",x"48",x"DF", -- 0x07B0
		x"94",x"FB",x"5D",x"4D",x"86",x"71",x"82",x"39", -- 0x07B8
		x"4B",x"B6",x"D4",x"86",x"57",x"2D",x"1C",x"F4", -- 0x07C0
		x"96",x"BF",x"C9",x"DF",x"19",x"7F",x"33",x"BC", -- 0x07C8
		x"6E",x"97",x"D8",x"FB",x"0F",x"22",x"DB",x"24", -- 0x07D0
		x"1E",x"39",x"F0",x"24",x"2A",x"F2",x"5D",x"76", -- 0x07D8
		x"29",x"B2",x"FC",x"81",x"DF",x"98",x"F5",x"F6", -- 0x07E0
		x"58",x"40",x"D6",x"72",x"BF",x"89",x"2F",x"AD", -- 0x07E8
		x"21",x"09",x"A9",x"AF",x"2B",x"06",x"53",x"C8", -- 0x07F0
		x"BE",x"44",x"ED",x"69",x"37",x"CA",x"DF",x"E0", -- 0x07F8
		x"7D",x"5C",x"62",x"DD",x"F5",x"58",x"54",x"CD", -- 0x0800
		x"18",x"AA",x"40",x"D7",x"34",x"EF",x"05",x"D4", -- 0x0808
		x"78",x"2F",x"84",x"23",x"35",x"D8",x"EB",x"73", -- 0x0810
		x"9C",x"59",x"DC",x"54",x"25",x"3C",x"35",x"22", -- 0x0818
		x"19",x"97",x"00",x"0F",x"6F",x"D3",x"5C",x"88", -- 0x0820
		x"7E",x"1D",x"DF",x"B2",x"0D",x"E5",x"87",x"05", -- 0x0828
		x"15",x"8C",x"28",x"C9",x"65",x"93",x"BC",x"81", -- 0x0830
		x"ED",x"9A",x"D5",x"13",x"56",x"0B",x"35",x"6F", -- 0x0838
		x"A2",x"B5",x"7E",x"92",x"89",x"DB",x"1B",x"88", -- 0x0840
		x"F8",x"7A",x"3B",x"85",x"DF",x"43",x"8A",x"74", -- 0x0848
		x"CF",x"32",x"3E",x"B4",x"C5",x"7B",x"36",x"B3", -- 0x0850
		x"16",x"0D",x"46",x"6C",x"97",x"FB",x"DC",x"BA", -- 0x0858
		x"B1",x"DA",x"4D",x"BA",x"36",x"E7",x"43",x"AE", -- 0x0860
		x"62",x"FE",x"34",x"43",x"C1",x"3E",x"B7",x"91", -- 0x0868
		x"70",x"76",x"C5",x"37",x"F1",x"7B",x"EA",x"87", -- 0x0870
		x"88",x"32",x"73",x"A0",x"AD",x"CF",x"5B",x"5F", -- 0x0878
		x"AB",x"A8",x"99",x"61",x"10",x"5D",x"11",x"F1", -- 0x0880
		x"DB",x"C4",x"35",x"9D",x"04",x"6D",x"AE",x"74", -- 0x0888
		x"63",x"74",x"2B",x"D4",x"EF",x"96",x"5C",x"F8", -- 0x0890
		x"48",x"CF",x"99",x"F5",x"20",x"74",x"D4",x"CB", -- 0x0898
		x"9C",x"6E",x"AC",x"AC",x"4B",x"BD",x"9E",x"27", -- 0x08A0
		x"83",x"54",x"C4",x"07",x"41",x"F2",x"7B",x"A4", -- 0x08A8
		x"67",x"27",x"79",x"D7",x"BD",x"55",x"50",x"06", -- 0x08B0
		x"A4",x"69",x"FB",x"C4",x"DD",x"D0",x"10",x"7A", -- 0x08B8
		x"BE",x"BD",x"A6",x"0B",x"FA",x"45",x"B1",x"7E", -- 0x08C0
		x"99",x"F6",x"85",x"DA",x"E9",x"81",x"FE",x"D1", -- 0x08C8
		x"A8",x"78",x"29",x"66",x"4D",x"79",x"EB",x"F2", -- 0x08D0
		x"62",x"67",x"37",x"BF",x"38",x"48",x"3A",x"76", -- 0x08D8
		x"06",x"60",x"01",x"01",x"A5",x"B3",x"00",x"BF", -- 0x08E0
		x"AA",x"05",x"9A",x"94",x"86",x"9A",x"E5",x"AE", -- 0x08E8
		x"92",x"0F",x"94",x"E0",x"08",x"80",x"53",x"6A", -- 0x08F0
		x"E7",x"8A",x"A9",x"9F",x"52",x"63",x"17",x"58", -- 0x08F8
		x"C3",x"18",x"D9",x"6A",x"4B",x"59",x"2A",x"F5", -- 0x0900
		x"5E",x"44",x"0B",x"65",x"5E",x"F0",x"14",x"F1", -- 0x0908
		x"80",x"29",x"52",x"88",x"A9",x"25",x"73",x"12", -- 0x0910
		x"2F",x"9C",x"31",x"82",x"01",x"48",x"5A",x"C4", -- 0x0918
		x"E0",x"B3",x"2F",x"2C",x"0D",x"D8",x"A2",x"EB", -- 0x0920
		x"1E",x"AD",x"51",x"FB",x"1E",x"E4",x"6D",x"9E", -- 0x0928
		x"8D",x"3F",x"A7",x"B7",x"64",x"9A",x"C9",x"94", -- 0x0930
		x"37",x"FA",x"17",x"38",x"C3",x"F0",x"7D",x"24", -- 0x0938
		x"A5",x"AC",x"50",x"B2",x"06",x"F2",x"1E",x"A3", -- 0x0940
		x"20",x"6F",x"9F",x"3F",x"D4",x"0E",x"5D",x"62", -- 0x0948
		x"4D",x"84",x"99",x"B2",x"1F",x"63",x"C6",x"D6", -- 0x0950
		x"DE",x"5D",x"0F",x"22",x"4E",x"8C",x"46",x"F3", -- 0x0958
		x"B9",x"16",x"27",x"3F",x"89",x"45",x"E2",x"29", -- 0x0960
		x"35",x"82",x"68",x"89",x"10",x"46",x"6B",x"5E", -- 0x0968
		x"CA",x"06",x"90",x"EA",x"E8",x"D6",x"C1",x"47", -- 0x0970
		x"B3",x"50",x"69",x"02",x"5D",x"2F",x"76",x"96", -- 0x0978
		x"C5",x"1D",x"D5",x"4F",x"62",x"B8",x"78",x"17", -- 0x0980
		x"BA",x"61",x"A0",x"CB",x"A7",x"8C",x"A9",x"F1", -- 0x0988
		x"92",x"B9",x"DC",x"7B",x"90",x"1E",x"C3",x"44", -- 0x0990
		x"EE",x"AC",x"C5",x"4C",x"DC",x"BB",x"62",x"A2", -- 0x0998
		x"D8",x"38",x"71",x"3C",x"70",x"69",x"D2",x"2B", -- 0x09A0
		x"CA",x"F3",x"76",x"F1",x"80",x"9F",x"E4",x"13", -- 0x09A8
		x"59",x"41",x"0E",x"69",x"DF",x"51",x"2D",x"CE", -- 0x09B0
		x"FE",x"F3",x"9A",x"5B",x"AF",x"FC",x"7D",x"89", -- 0x09B8
		x"B4",x"EE",x"45",x"25",x"D7",x"97",x"CF",x"A3", -- 0x09C0
		x"8B",x"C6",x"15",x"0C",x"66",x"F9",x"9E",x"40", -- 0x09C8
		x"3C",x"AD",x"29",x"1C",x"7E",x"57",x"6A",x"7D", -- 0x09D0
		x"CA",x"05",x"58",x"7A",x"81",x"D5",x"83",x"36", -- 0x09D8
		x"44",x"48",x"5B",x"1D",x"E0",x"2B",x"40",x"EB", -- 0x09E0
		x"71",x"55",x"F8",x"D8",x"CF",x"97",x"98",x"0C", -- 0x09E8
		x"C4",x"C1",x"A7",x"44",x"19",x"12",x"41",x"E3", -- 0x09F0
		x"96",x"9A",x"DE",x"18",x"EF",x"E1",x"4E",x"B4", -- 0x09F8
		x"AA",x"29",x"51",x"8B",x"D3",x"91",x"F6",x"46", -- 0x0A00
		x"66",x"EF",x"9E",x"36",x"08",x"37",x"C1",x"CC", -- 0x0A08
		x"78",x"69",x"90",x"92",x"FA",x"D2",x"F5",x"11", -- 0x0A10
		x"EC",x"54",x"29",x"DC",x"37",x"F6",x"11",x"E1", -- 0x0A18
		x"9F",x"62",x"EC",x"74",x"F3",x"E3",x"3A",x"DA", -- 0x0A20
		x"54",x"D8",x"90",x"5C",x"8F",x"53",x"A8",x"08", -- 0x0A28
		x"3C",x"3A",x"1A",x"B7",x"8C",x"11",x"C8",x"79", -- 0x0A30
		x"E4",x"72",x"D5",x"1C",x"69",x"E7",x"7D",x"89", -- 0x0A38
		x"4A",x"6A",x"FD",x"BE",x"CE",x"38",x"19",x"23", -- 0x0A40
		x"90",x"A9",x"FE",x"20",x"FC",x"A7",x"28",x"B9", -- 0x0A48
		x"E1",x"C2",x"71",x"6E",x"53",x"3A",x"67",x"38", -- 0x0A50
		x"AC",x"3E",x"D4",x"96",x"A5",x"52",x"20",x"6F", -- 0x0A58
		x"3D",x"1E",x"AD",x"0C",x"D5",x"C6",x"AE",x"E5", -- 0x0A60
		x"F0",x"AD",x"06",x"ED",x"55",x"AD",x"27",x"B7", -- 0x0A68
		x"70",x"98",x"A5",x"C3",x"D3",x"8D",x"FC",x"00", -- 0x0A70
		x"4B",x"51",x"96",x"F0",x"A3",x"B6",x"DF",x"E0", -- 0x0A78
		x"54",x"8E",x"6C",x"A9",x"D4",x"1B",x"8F",x"C5", -- 0x0A80
		x"48",x"95",x"34",x"1E",x"C3",x"5B",x"D5",x"34", -- 0x0A88
		x"F4",x"FA",x"78",x"48",x"88",x"F4",x"48",x"D3", -- 0x0A90
		x"46",x"DF",x"44",x"E9",x"16",x"25",x"4B",x"6B", -- 0x0A98
		x"33",x"B7",x"15",x"08",x"53",x"A5",x"4E",x"1B", -- 0x0AA0
		x"BA",x"82",x"39",x"7E",x"5D",x"8E",x"B3",x"D1", -- 0x0AA8
		x"8A",x"2C",x"1A",x"92",x"21",x"E2",x"E6",x"E6", -- 0x0AB0
		x"C2",x"2B",x"D0",x"D8",x"50",x"9B",x"C3",x"83", -- 0x0AB8
		x"54",x"D9",x"0C",x"27",x"FE",x"5A",x"C1",x"B9", -- 0x0AC0
		x"DC",x"FB",x"39",x"3A",x"8A",x"6C",x"0D",x"94", -- 0x0AC8
		x"18",x"A6",x"A7",x"B8",x"89",x"8E",x"9F",x"CB", -- 0x0AD0
		x"B9",x"70",x"25",x"8A",x"0D",x"E8",x"0E",x"E0", -- 0x0AD8
		x"42",x"1A",x"87",x"41",x"74",x"49",x"FB",x"D0", -- 0x0AE0
		x"C4",x"B4",x"8B",x"CF",x"21",x"18",x"64",x"39", -- 0x0AE8
		x"BE",x"0C",x"F1",x"C8",x"1A",x"91",x"94",x"D4", -- 0x0AF0
		x"81",x"39",x"5F",x"0E",x"23",x"EC",x"6E",x"65", -- 0x0AF8
		x"08",x"75",x"A7",x"FB",x"BF",x"23",x"4D",x"04", -- 0x0B00
		x"D7",x"D8",x"D3",x"F8",x"70",x"B8",x"B1",x"AE", -- 0x0B08
		x"44",x"23",x"77",x"5F",x"B4",x"8C",x"34",x"B5", -- 0x0B10
		x"C5",x"13",x"C4",x"68",x"00",x"B2",x"CE",x"87", -- 0x0B18
		x"29",x"F5",x"04",x"68",x"19",x"51",x"6C",x"70", -- 0x0B20
		x"A9",x"41",x"E8",x"99",x"F9",x"9A",x"48",x"BD", -- 0x0B28
		x"BD",x"40",x"1D",x"F1",x"CC",x"D0",x"27",x"12", -- 0x0B30
		x"E3",x"6B",x"7B",x"64",x"1F",x"C9",x"EB",x"48", -- 0x0B38
		x"3F",x"6F",x"B0",x"D7",x"40",x"9C",x"48",x"69", -- 0x0B40
		x"DD",x"31",x"03",x"57",x"4B",x"4C",x"16",x"88", -- 0x0B48
		x"8C",x"B2",x"F9",x"D8",x"84",x"21",x"EA",x"E7", -- 0x0B50
		x"8D",x"E5",x"4C",x"AC",x"2F",x"B8",x"74",x"6E", -- 0x0B58
		x"28",x"A4",x"46",x"E8",x"41",x"0E",x"52",x"20", -- 0x0B60
		x"3F",x"56",x"F6",x"0A",x"A2",x"8C",x"92",x"AE", -- 0x0B68
		x"40",x"8C",x"07",x"44",x"2E",x"F1",x"2C",x"BB", -- 0x0B70
		x"58",x"F8",x"68",x"87",x"31",x"5C",x"76",x"D8", -- 0x0B78
		x"01",x"BC",x"C1",x"42",x"CB",x"15",x"62",x"8A", -- 0x0B80
		x"6B",x"D9",x"15",x"8D",x"66",x"27",x"3C",x"26", -- 0x0B88
		x"34",x"43",x"6A",x"62",x"B4",x"17",x"1E",x"8C", -- 0x0B90
		x"8F",x"06",x"94",x"C0",x"62",x"0B",x"99",x"E2", -- 0x0B98
		x"47",x"5C",x"25",x"92",x"71",x"08",x"1E",x"5C", -- 0x0BA0
		x"E1",x"B2",x"E9",x"C7",x"D9",x"A5",x"EE",x"0E", -- 0x0BA8
		x"68",x"59",x"EF",x"9C",x"EF",x"0E",x"A9",x"7F", -- 0x0BB0
		x"93",x"3E",x"40",x"75",x"49",x"DA",x"58",x"10", -- 0x0BB8
		x"B6",x"7E",x"A3",x"A7",x"06",x"41",x"83",x"E7", -- 0x0BC0
		x"F3",x"6D",x"AF",x"4D",x"92",x"1E",x"DB",x"7A", -- 0x0BC8
		x"F7",x"CB",x"17",x"E7",x"DA",x"C0",x"68",x"ED", -- 0x0BD0
		x"7E",x"A8",x"E3",x"47",x"03",x"3C",x"58",x"39", -- 0x0BD8
		x"3A",x"7B",x"60",x"40",x"BC",x"E3",x"A7",x"30", -- 0x0BE0
		x"D0",x"D7",x"7D",x"63",x"F5",x"59",x"5D",x"ED", -- 0x0BE8
		x"26",x"75",x"D6",x"80",x"B5",x"BE",x"ED",x"B4", -- 0x0BF0
		x"E6",x"D1",x"FB",x"6A",x"8E",x"54",x"A3",x"C8", -- 0x0BF8
		x"4F",x"05",x"89",x"0C",x"E8",x"31",x"BB",x"3A", -- 0x0C00
		x"09",x"B9",x"9D",x"7F",x"13",x"FB",x"6D",x"B8", -- 0x0C08
		x"F0",x"C3",x"B8",x"26",x"82",x"27",x"DA",x"6A", -- 0x0C10
		x"F8",x"57",x"D4",x"07",x"AB",x"F7",x"D0",x"7B", -- 0x0C18
		x"7C",x"5A",x"87",x"E5",x"0B",x"C3",x"20",x"15", -- 0x0C20
		x"7D",x"3D",x"94",x"10",x"B8",x"81",x"49",x"29", -- 0x0C28
		x"46",x"81",x"50",x"48",x"A8",x"AA",x"32",x"22", -- 0x0C30
		x"02",x"86",x"29",x"2E",x"7F",x"79",x"A9",x"FB", -- 0x0C38
		x"D3",x"B0",x"61",x"DF",x"74",x"81",x"74",x"71", -- 0x0C40
		x"BF",x"88",x"02",x"78",x"0A",x"4B",x"A2",x"CF", -- 0x0C48
		x"CC",x"72",x"19",x"F5",x"1D",x"CA",x"18",x"9F", -- 0x0C50
		x"52",x"C0",x"CD",x"D1",x"3B",x"F6",x"4D",x"8E", -- 0x0C58
		x"A7",x"AF",x"ED",x"9C",x"B0",x"62",x"8D",x"70", -- 0x0C60
		x"6A",x"8F",x"69",x"75",x"DA",x"8B",x"C4",x"28", -- 0x0C68
		x"FD",x"DD",x"9D",x"9A",x"A9",x"35",x"B9",x"7B", -- 0x0C70
		x"F5",x"07",x"4D",x"B0",x"FD",x"1A",x"40",x"26", -- 0x0C78
		x"49",x"2E",x"42",x"FA",x"11",x"CF",x"6B",x"7B", -- 0x0C80
		x"60",x"54",x"70",x"BA",x"DF",x"36",x"62",x"5D", -- 0x0C88
		x"93",x"00",x"78",x"BC",x"35",x"B1",x"38",x"AB", -- 0x0C90
		x"B9",x"05",x"5C",x"B7",x"20",x"1C",x"5D",x"E8", -- 0x0C98
		x"CA",x"9F",x"E3",x"5B",x"EF",x"CF",x"56",x"50", -- 0x0CA0
		x"24",x"C7",x"8A",x"84",x"7D",x"6D",x"61",x"11", -- 0x0CA8
		x"6D",x"59",x"CE",x"23",x"0C",x"86",x"4E",x"45", -- 0x0CB0
		x"8C",x"AA",x"7C",x"2C",x"47",x"DA",x"15",x"12", -- 0x0CB8
		x"F9",x"79",x"EC",x"E9",x"49",x"43",x"B9",x"EC", -- 0x0CC0
		x"0B",x"45",x"F0",x"08",x"B2",x"53",x"1A",x"9F", -- 0x0CC8
		x"2C",x"68",x"C2",x"B7",x"EE",x"90",x"FC",x"FA", -- 0x0CD0
		x"BB",x"7A",x"A6",x"03",x"D4",x"3C",x"94",x"CE", -- 0x0CD8
		x"B5",x"81",x"B9",x"FE",x"44",x"F2",x"6B",x"50", -- 0x0CE0
		x"38",x"5D",x"D7",x"6A",x"B0",x"F1",x"0B",x"5C", -- 0x0CE8
		x"D9",x"4D",x"15",x"C9",x"DE",x"91",x"44",x"9A", -- 0x0CF0
		x"0C",x"EB",x"1D",x"60",x"28",x"31",x"AF",x"DD", -- 0x0CF8
		x"B2",x"E8",x"5C",x"F6",x"DB",x"C7",x"C6",x"15", -- 0x0D00
		x"25",x"9F",x"FE",x"55",x"11",x"0A",x"32",x"EB", -- 0x0D08
		x"D7",x"47",x"35",x"36",x"D8",x"79",x"50",x"65", -- 0x0D10
		x"E4",x"6D",x"45",x"8C",x"1E",x"F4",x"6A",x"D0", -- 0x0D18
		x"DD",x"46",x"47",x"BA",x"0F",x"8E",x"4F",x"B3", -- 0x0D20
		x"AD",x"4E",x"89",x"BE",x"D8",x"BB",x"2A",x"B0", -- 0x0D28
		x"82",x"5F",x"66",x"DA",x"59",x"B6",x"BF",x"3E", -- 0x0D30
		x"A3",x"06",x"CB",x"C1",x"FA",x"B5",x"12",x"59", -- 0x0D38
		x"FC",x"D8",x"14",x"8B",x"67",x"63",x"BE",x"15", -- 0x0D40
		x"31",x"C7",x"54",x"0A",x"83",x"7E",x"3A",x"06", -- 0x0D48
		x"DE",x"A0",x"E1",x"38",x"D6",x"21",x"F5",x"F9", -- 0x0D50
		x"27",x"C1",x"BB",x"23",x"F7",x"4D",x"FB",x"74", -- 0x0D58
		x"27",x"10",x"7F",x"0E",x"F2",x"BD",x"24",x"24", -- 0x0D60
		x"86",x"F7",x"AE",x"0A",x"76",x"E8",x"90",x"D4", -- 0x0D68
		x"8A",x"F1",x"0D",x"E0",x"13",x"83",x"DB",x"3B", -- 0x0D70
		x"C4",x"17",x"DD",x"BC",x"65",x"59",x"31",x"0C", -- 0x0D78
		x"69",x"30",x"1A",x"DB",x"EE",x"BD",x"00",x"75", -- 0x0D80
		x"B5",x"AE",x"FE",x"AC",x"18",x"0F",x"81",x"22", -- 0x0D88
		x"01",x"0F",x"03",x"94",x"92",x"DE",x"4F",x"57", -- 0x0D90
		x"F6",x"AC",x"15",x"DB",x"06",x"C5",x"E7",x"EE", -- 0x0D98
		x"76",x"02",x"CA",x"65",x"40",x"4A",x"5A",x"F5", -- 0x0DA0
		x"79",x"59",x"A2",x"91",x"69",x"A4",x"B3",x"E9", -- 0x0DA8
		x"B3",x"B6",x"FD",x"46",x"16",x"4D",x"9D",x"0D", -- 0x0DB0
		x"79",x"32",x"E8",x"7F",x"78",x"D0",x"6E",x"6E", -- 0x0DB8
		x"52",x"B8",x"D3",x"92",x"04",x"AD",x"09",x"7D", -- 0x0DC0
		x"07",x"2B",x"8E",x"EF",x"CF",x"42",x"5A",x"83", -- 0x0DC8
		x"78",x"D7",x"49",x"8E",x"26",x"67",x"1B",x"9F", -- 0x0DD0
		x"19",x"04",x"9F",x"11",x"54",x"8D",x"7F",x"27", -- 0x0DD8
		x"47",x"53",x"39",x"CA",x"80",x"42",x"C7",x"08", -- 0x0DE0
		x"ED",x"D5",x"F7",x"BD",x"18",x"D1",x"C1",x"10", -- 0x0DE8
		x"AA",x"0B",x"1F",x"50",x"F1",x"3A",x"6F",x"0C", -- 0x0DF0
		x"BE",x"8E",x"1D",x"13",x"1D",x"9D",x"B9",x"E3", -- 0x0DF8
		x"70",x"F3",x"AE",x"F1",x"36",x"F5",x"F9",x"24", -- 0x0E00
		x"CB",x"71",x"62",x"63",x"C3",x"24",x"73",x"ED", -- 0x0E08
		x"AE",x"12",x"3E",x"A1",x"4D",x"2D",x"2D",x"0C", -- 0x0E10
		x"BC",x"4A",x"9E",x"D9",x"67",x"59",x"BD",x"58", -- 0x0E18
		x"4D",x"EB",x"4A",x"03",x"61",x"C3",x"A7",x"2D", -- 0x0E20
		x"B4",x"0A",x"90",x"78",x"AD",x"83",x"66",x"DB", -- 0x0E28
		x"16",x"24",x"7D",x"63",x"52",x"2A",x"EE",x"0F", -- 0x0E30
		x"F4",x"8D",x"68",x"5C",x"66",x"A5",x"B4",x"B3", -- 0x0E38
		x"11",x"7E",x"37",x"72",x"C1",x"DE",x"9F",x"77", -- 0x0E40
		x"E8",x"AF",x"6F",x"96",x"B2",x"D6",x"F1",x"C8", -- 0x0E48
		x"7A",x"70",x"AB",x"CC",x"1A",x"9A",x"5B",x"0F", -- 0x0E50
		x"A8",x"C3",x"6C",x"8E",x"E8",x"A0",x"43",x"F9", -- 0x0E58
		x"9F",x"7A",x"6C",x"61",x"D8",x"8B",x"58",x"C1", -- 0x0E60
		x"BA",x"C8",x"D7",x"6E",x"9F",x"C9",x"B6",x"99", -- 0x0E68
		x"B9",x"E2",x"67",x"D4",x"FC",x"42",x"E3",x"A5", -- 0x0E70
		x"86",x"CF",x"35",x"6F",x"F0",x"F7",x"6A",x"10", -- 0x0E78
		x"F1",x"56",x"71",x"CA",x"E2",x"CA",x"0C",x"9D", -- 0x0E80
		x"93",x"E3",x"8B",x"B2",x"2D",x"C2",x"4C",x"E7", -- 0x0E88
		x"A5",x"33",x"3C",x"A2",x"F5",x"9F",x"C8",x"7C", -- 0x0E90
		x"EF",x"7D",x"EB",x"60",x"F4",x"D5",x"70",x"66", -- 0x0E98
		x"2D",x"61",x"B0",x"8F",x"2C",x"BC",x"2D",x"3F", -- 0x0EA0
		x"20",x"39",x"71",x"CC",x"FB",x"3E",x"B4",x"21", -- 0x0EA8
		x"71",x"70",x"43",x"67",x"90",x"8B",x"63",x"80", -- 0x0EB0
		x"88",x"CF",x"E0",x"7D",x"A5",x"D0",x"63",x"52", -- 0x0EB8
		x"32",x"14",x"E1",x"DE",x"50",x"10",x"1E",x"70", -- 0x0EC0
		x"C8",x"90",x"3E",x"44",x"CE",x"72",x"65",x"BF", -- 0x0EC8
		x"63",x"28",x"A7",x"F3",x"B4",x"0B",x"74",x"3D", -- 0x0ED0
		x"DA",x"D4",x"3B",x"01",x"A5",x"9E",x"53",x"57", -- 0x0ED8
		x"B3",x"36",x"36",x"04",x"C5",x"55",x"F4",x"8E", -- 0x0EE0
		x"65",x"B2",x"D2",x"B3",x"25",x"B7",x"F2",x"88", -- 0x0EE8
		x"DF",x"9A",x"FB",x"14",x"26",x"EF",x"52",x"80", -- 0x0EF0
		x"C4",x"8D",x"81",x"E9",x"AB",x"55",x"42",x"DE", -- 0x0EF8
		x"8B",x"78",x"E3",x"D0",x"4D",x"58",x"DE",x"32", -- 0x0F00
		x"0B",x"31",x"65",x"AF",x"E8",x"59",x"B8",x"48", -- 0x0F08
		x"73",x"B4",x"5D",x"19",x"A5",x"2F",x"1A",x"E9", -- 0x0F10
		x"3C",x"9B",x"D4",x"E7",x"70",x"96",x"C7",x"7B", -- 0x0F18
		x"8E",x"2B",x"4C",x"5C",x"03",x"2B",x"8E",x"0E", -- 0x0F20
		x"5C",x"74",x"3D",x"C4",x"4D",x"F5",x"0E",x"C0", -- 0x0F28
		x"2B",x"EA",x"5A",x"D0",x"99",x"74",x"BA",x"D5", -- 0x0F30
		x"8F",x"0F",x"3D",x"01",x"A5",x"05",x"7C",x"B4", -- 0x0F38
		x"AF",x"49",x"11",x"B2",x"74",x"1F",x"40",x"D1", -- 0x0F40
		x"93",x"7E",x"96",x"60",x"F3",x"24",x"22",x"1F", -- 0x0F48
		x"8E",x"FB",x"EF",x"28",x"70",x"2B",x"FD",x"7F", -- 0x0F50
		x"B9",x"3C",x"00",x"DF",x"C0",x"7D",x"94",x"F0", -- 0x0F58
		x"C6",x"25",x"23",x"BA",x"44",x"64",x"8C",x"58", -- 0x0F60
		x"62",x"A3",x"B8",x"D5",x"47",x"5A",x"F5",x"D6", -- 0x0F68
		x"D5",x"65",x"FE",x"C5",x"10",x"7D",x"46",x"CA", -- 0x0F70
		x"39",x"46",x"AA",x"F9",x"43",x"3F",x"6A",x"0A", -- 0x0F78
		x"E3",x"8E",x"C5",x"28",x"72",x"D1",x"00",x"D4", -- 0x0F80
		x"F4",x"39",x"AA",x"3D",x"93",x"20",x"93",x"6A", -- 0x0F88
		x"86",x"92",x"30",x"16",x"10",x"F5",x"E0",x"C8", -- 0x0F90
		x"3D",x"8B",x"C3",x"80",x"4A",x"AD",x"0B",x"2E", -- 0x0F98
		x"3C",x"50",x"D6",x"AE",x"22",x"56",x"03",x"97", -- 0x0FA0
		x"8F",x"2E",x"D4",x"A3",x"CD",x"E7",x"8D",x"D3", -- 0x0FA8
		x"7A",x"3D",x"EA",x"0B",x"34",x"CB",x"D3",x"71", -- 0x0FB0
		x"D7",x"17",x"71",x"A1",x"C5",x"7C",x"50",x"81", -- 0x0FB8
		x"4C",x"A6",x"B0",x"6F",x"FC",x"B3",x"86",x"0D", -- 0x0FC0
		x"61",x"DA",x"B0",x"30",x"C2",x"3E",x"83",x"3D", -- 0x0FC8
		x"7B",x"6E",x"C7",x"2F",x"BA",x"1C",x"A0",x"92", -- 0x0FD0
		x"B2",x"92",x"B3",x"F7",x"8E",x"04",x"7A",x"DB", -- 0x0FD8
		x"AA",x"2B",x"CA",x"28",x"5E",x"51",x"35",x"40", -- 0x0FE0
		x"2C",x"65",x"EF",x"EE",x"23",x"73",x"AB",x"9E", -- 0x0FE8
		x"62",x"F3",x"4E",x"1D",x"10",x"EE",x"2F",x"42", -- 0x0FF0
		x"01",x"E2",x"3B",x"90",x"67",x"B5",x"6C",x"12", -- 0x0FF8
		x"60",x"37",x"B9",x"3E",x"88",x"6E",x"FD",x"34", -- 0x1000
		x"D3",x"ED",x"23",x"F6",x"E1",x"4E",x"16",x"44", -- 0x1008
		x"42",x"64",x"E0",x"D1",x"D2",x"10",x"15",x"D4", -- 0x1010
		x"F2",x"50",x"E4",x"5A",x"85",x"51",x"EC",x"65", -- 0x1018
		x"88",x"26",x"23",x"90",x"95",x"22",x"C4",x"E8", -- 0x1020
		x"8F",x"67",x"E0",x"71",x"B5",x"76",x"35",x"F8", -- 0x1028
		x"5A",x"16",x"CA",x"AC",x"A5",x"5F",x"01",x"19", -- 0x1030
		x"2F",x"E5",x"73",x"34",x"37",x"DF",x"99",x"3F", -- 0x1038
		x"07",x"3D",x"CF",x"1C",x"5F",x"14",x"05",x"6E", -- 0x1040
		x"7B",x"65",x"60",x"32",x"DB",x"95",x"AA",x"B5", -- 0x1048
		x"2C",x"F4",x"63",x"D1",x"55",x"64",x"EA",x"04", -- 0x1050
		x"CA",x"DE",x"39",x"02",x"3E",x"D2",x"42",x"45", -- 0x1058
		x"10",x"91",x"E0",x"EE",x"26",x"E6",x"5E",x"A1", -- 0x1060
		x"4C",x"BE",x"53",x"A8",x"D3",x"FD",x"DD",x"00", -- 0x1068
		x"F3",x"41",x"52",x"C8",x"26",x"3D",x"CC",x"F0", -- 0x1070
		x"9B",x"06",x"72",x"DA",x"59",x"34",x"9F",x"E8", -- 0x1078
		x"C6",x"81",x"58",x"EC",x"E7",x"B6",x"0E",x"34", -- 0x1080
		x"F4",x"62",x"5C",x"C8",x"DF",x"3B",x"49",x"53", -- 0x1088
		x"FB",x"9B",x"1C",x"22",x"58",x"69",x"92",x"74", -- 0x1090
		x"EE",x"06",x"4F",x"C7",x"3A",x"6E",x"B1",x"80", -- 0x1098
		x"EF",x"0A",x"EC",x"57",x"40",x"7B",x"8C",x"35", -- 0x10A0
		x"DD",x"68",x"7D",x"BD",x"A3",x"46",x"91",x"20", -- 0x10A8
		x"E1",x"2D",x"C1",x"BA",x"96",x"55",x"2F",x"06", -- 0x10B0
		x"DA",x"FD",x"CD",x"94",x"6C",x"FE",x"95",x"DC", -- 0x10B8
		x"88",x"82",x"B3",x"C8",x"FD",x"BF",x"7D",x"5B", -- 0x10C0
		x"29",x"7B",x"99",x"4C",x"C1",x"2B",x"6C",x"24", -- 0x10C8
		x"58",x"2F",x"5E",x"6F",x"04",x"8D",x"75",x"DE", -- 0x10D0
		x"0B",x"C2",x"F2",x"F6",x"C2",x"88",x"53",x"CA", -- 0x10D8
		x"8B",x"08",x"94",x"09",x"C7",x"91",x"65",x"70", -- 0x10E0
		x"8C",x"7E",x"BD",x"4F",x"A9",x"2A",x"F2",x"81", -- 0x10E8
		x"59",x"51",x"F0",x"5D",x"5E",x"E5",x"BB",x"69", -- 0x10F0
		x"29",x"AF",x"DF",x"6B",x"38",x"B3",x"36",x"43", -- 0x10F8
		x"BB",x"4A",x"4D",x"03",x"5C",x"32",x"74",x"E8", -- 0x1100
		x"B0",x"32",x"B7",x"5A",x"DB",x"AA",x"5B",x"B5", -- 0x1108
		x"FB",x"CC",x"92",x"5A",x"32",x"CE",x"43",x"5B", -- 0x1110
		x"7E",x"24",x"46",x"36",x"D7",x"7D",x"7A",x"13", -- 0x1118
		x"47",x"47",x"16",x"A3",x"79",x"0A",x"8D",x"2A", -- 0x1120
		x"BB",x"45",x"04",x"98",x"70",x"DE",x"CD",x"6C", -- 0x1128
		x"AB",x"DF",x"C7",x"DE",x"AE",x"0B",x"B9",x"AC", -- 0x1130
		x"AE",x"01",x"E3",x"06",x"FD",x"DD",x"19",x"45", -- 0x1138
		x"A4",x"AF",x"69",x"1E",x"B9",x"F6",x"C7",x"F5", -- 0x1140
		x"BB",x"CB",x"0E",x"2C",x"AA",x"DB",x"19",x"D6", -- 0x1148
		x"BB",x"60",x"35",x"EA",x"EA",x"EE",x"97",x"9A", -- 0x1150
		x"6F",x"7B",x"A0",x"EC",x"D8",x"3A",x"33",x"7D", -- 0x1158
		x"E9",x"9C",x"9B",x"23",x"13",x"63",x"19",x"4E", -- 0x1160
		x"AE",x"27",x"FA",x"D9",x"82",x"14",x"B0",x"BE", -- 0x1168
		x"74",x"E5",x"A9",x"5F",x"54",x"41",x"79",x"44", -- 0x1170
		x"3D",x"9A",x"31",x"16",x"D4",x"64",x"14",x"3E", -- 0x1178
		x"80",x"2F",x"61",x"13",x"13",x"FA",x"62",x"C1", -- 0x1180
		x"A1",x"DC",x"1B",x"25",x"70",x"CB",x"E3",x"64", -- 0x1188
		x"31",x"0D",x"43",x"86",x"4E",x"BD",x"CA",x"8B", -- 0x1190
		x"58",x"FB",x"22",x"AC",x"E0",x"36",x"6A",x"E0", -- 0x1198
		x"65",x"CB",x"F4",x"F7",x"46",x"D6",x"BA",x"E8", -- 0x11A0
		x"B3",x"D5",x"8D",x"A3",x"22",x"F0",x"08",x"53", -- 0x11A8
		x"FD",x"4B",x"59",x"4C",x"09",x"24",x"58",x"E0", -- 0x11B0
		x"A0",x"7A",x"0D",x"81",x"30",x"77",x"E1",x"15", -- 0x11B8
		x"C3",x"D6",x"0E",x"0A",x"AD",x"48",x"72",x"E0", -- 0x11C0
		x"9D",x"7F",x"84",x"BF",x"70",x"8C",x"93",x"6E", -- 0x11C8
		x"58",x"EC",x"3B",x"E0",x"91",x"93",x"C2",x"32", -- 0x11D0
		x"8D",x"4F",x"33",x"BD",x"C7",x"15",x"D2",x"0B", -- 0x11D8
		x"6C",x"E0",x"94",x"99",x"A8",x"08",x"7B",x"47", -- 0x11E0
		x"87",x"7F",x"86",x"78",x"8C",x"1A",x"E6",x"E4", -- 0x11E8
		x"87",x"22",x"C5",x"19",x"35",x"08",x"CA",x"C2", -- 0x11F0
		x"58",x"7D",x"80",x"9F",x"12",x"D3",x"AA",x"7E", -- 0x11F8
		x"34",x"3F",x"19",x"DD",x"C6",x"14",x"A4",x"CE", -- 0x1200
		x"13",x"2B",x"47",x"9F",x"C5",x"AD",x"04",x"CC", -- 0x1208
		x"D0",x"CA",x"E5",x"85",x"52",x"30",x"49",x"2A", -- 0x1210
		x"2D",x"C9",x"C9",x"3F",x"1D",x"F3",x"3E",x"52", -- 0x1218
		x"34",x"D6",x"30",x"FA",x"EA",x"D4",x"49",x"7D", -- 0x1220
		x"7F",x"90",x"9D",x"45",x"3F",x"A1",x"12",x"8F", -- 0x1228
		x"EB",x"77",x"15",x"3F",x"27",x"5E",x"69",x"54", -- 0x1230
		x"A8",x"34",x"14",x"C5",x"28",x"52",x"18",x"DB", -- 0x1238
		x"29",x"C7",x"57",x"93",x"1C",x"A0",x"11",x"9C", -- 0x1240
		x"B1",x"AE",x"61",x"F0",x"D0",x"F3",x"80",x"BC", -- 0x1248
		x"EA",x"15",x"FB",x"13",x"F3",x"66",x"E6",x"9C", -- 0x1250
		x"1A",x"7A",x"E1",x"C1",x"CC",x"7A",x"1E",x"75", -- 0x1258
		x"42",x"75",x"09",x"5F",x"95",x"9A",x"7B",x"47", -- 0x1260
		x"C8",x"DC",x"38",x"99",x"50",x"38",x"57",x"3C", -- 0x1268
		x"CD",x"D2",x"CE",x"C1",x"B8",x"35",x"DD",x"D2", -- 0x1270
		x"B0",x"BF",x"15",x"7D",x"B9",x"33",x"F3",x"FC", -- 0x1278
		x"28",x"7C",x"DB",x"BD",x"17",x"57",x"06",x"60", -- 0x1280
		x"B3",x"BD",x"F9",x"05",x"76",x"D0",x"C0",x"C3", -- 0x1288
		x"A4",x"8F",x"85",x"5D",x"C4",x"63",x"B0",x"75", -- 0x1290
		x"A2",x"C5",x"73",x"5D",x"78",x"67",x"D9",x"A0", -- 0x1298
		x"63",x"35",x"5E",x"FA",x"0C",x"E3",x"5B",x"BF", -- 0x12A0
		x"22",x"D4",x"44",x"18",x"26",x"05",x"DB",x"CA", -- 0x12A8
		x"94",x"61",x"A7",x"D9",x"44",x"D7",x"CE",x"66", -- 0x12B0
		x"1D",x"42",x"43",x"95",x"29",x"1D",x"B5",x"8D", -- 0x12B8
		x"D1",x"94",x"88",x"DD",x"F7",x"63",x"9E",x"1A", -- 0x12C0
		x"B7",x"62",x"32",x"DD",x"68",x"0E",x"28",x"7C", -- 0x12C8
		x"EE",x"D0",x"D5",x"33",x"28",x"A5",x"1A",x"C5", -- 0x12D0
		x"E7",x"5D",x"5B",x"91",x"FA",x"91",x"9E",x"CC", -- 0x12D8
		x"26",x"A6",x"AB",x"9D",x"0A",x"C9",x"B8",x"C1", -- 0x12E0
		x"2C",x"EA",x"A0",x"14",x"79",x"C8",x"11",x"68", -- 0x12E8
		x"19",x"E6",x"1C",x"C1",x"0C",x"36",x"87",x"74", -- 0x12F0
		x"13",x"62",x"06",x"0E",x"F3",x"A4",x"DB",x"99", -- 0x12F8
		x"4B",x"07",x"38",x"D4",x"50",x"70",x"16",x"FB", -- 0x1300
		x"DA",x"B6",x"11",x"54",x"00",x"A1",x"3D",x"98", -- 0x1308
		x"08",x"59",x"D9",x"15",x"0F",x"61",x"89",x"22", -- 0x1310
		x"C4",x"8F",x"31",x"38",x"B3",x"8C",x"52",x"7E", -- 0x1318
		x"13",x"0A",x"53",x"63",x"7A",x"69",x"5F",x"55", -- 0x1320
		x"A0",x"EF",x"2A",x"20",x"11",x"67",x"38",x"1A", -- 0x1328
		x"40",x"13",x"2F",x"CE",x"74",x"B8",x"F0",x"B8", -- 0x1330
		x"C7",x"A1",x"71",x"FA",x"AD",x"C3",x"79",x"40", -- 0x1338
		x"CD",x"CC",x"A3",x"C7",x"B5",x"83",x"9C",x"D5", -- 0x1340
		x"F2",x"46",x"F5",x"05",x"2D",x"2F",x"9E",x"6D", -- 0x1348
		x"42",x"CD",x"3C",x"36",x"06",x"AD",x"EF",x"4D", -- 0x1350
		x"CE",x"61",x"48",x"7D",x"A4",x"C1",x"BD",x"F1", -- 0x1358
		x"0E",x"E1",x"B9",x"C3",x"E4",x"D5",x"1A",x"57", -- 0x1360
		x"1D",x"10",x"DB",x"4A",x"BE",x"7A",x"B8",x"01", -- 0x1368
		x"48",x"74",x"B7",x"CD",x"A1",x"A7",x"1B",x"71", -- 0x1370
		x"88",x"63",x"6E",x"2D",x"A4",x"AB",x"1F",x"B2", -- 0x1378
		x"8D",x"58",x"F6",x"F1",x"2E",x"11",x"4A",x"4B", -- 0x1380
		x"A0",x"26",x"96",x"60",x"A1",x"CE",x"E0",x"69", -- 0x1388
		x"C2",x"98",x"38",x"65",x"BF",x"D2",x"56",x"48", -- 0x1390
		x"B6",x"C4",x"75",x"5B",x"70",x"14",x"8E",x"7E", -- 0x1398
		x"6C",x"85",x"70",x"9B",x"16",x"BA",x"66",x"B6", -- 0x13A0
		x"61",x"FC",x"96",x"82",x"4B",x"78",x"EB",x"0F", -- 0x13A8
		x"11",x"A3",x"74",x"D1",x"77",x"4A",x"99",x"2E", -- 0x13B0
		x"0F",x"10",x"09",x"FE",x"A3",x"97",x"7D",x"11", -- 0x13B8
		x"9C",x"EE",x"2C",x"B2",x"29",x"92",x"E9",x"0A", -- 0x13C0
		x"10",x"80",x"8C",x"5B",x"F8",x"F8",x"6A",x"8A", -- 0x13C8
		x"9C",x"5E",x"DB",x"93",x"A8",x"75",x"41",x"37", -- 0x13D0
		x"05",x"CA",x"37",x"A9",x"62",x"B4",x"3A",x"7F", -- 0x13D8
		x"A3",x"66",x"32",x"4D",x"78",x"9B",x"57",x"88", -- 0x13E0
		x"1D",x"64",x"E4",x"95",x"5D",x"4F",x"9F",x"79", -- 0x13E8
		x"2E",x"7B",x"8D",x"D6",x"F1",x"CE",x"0F",x"76", -- 0x13F0
		x"99",x"46",x"20",x"7C",x"FA",x"D9",x"FB",x"1F", -- 0x13F8
		x"40",x"AD",x"EB",x"B9",x"4A",x"C2",x"C1",x"E6", -- 0x1400
		x"27",x"A6",x"FB",x"04",x"76",x"9C",x"7E",x"A4", -- 0x1408
		x"97",x"0C",x"7B",x"09",x"5A",x"0A",x"80",x"74", -- 0x1410
		x"50",x"20",x"F0",x"CB",x"FA",x"6C",x"EA",x"BA", -- 0x1418
		x"1A",x"56",x"F3",x"E3",x"19",x"B6",x"4A",x"C0", -- 0x1420
		x"DC",x"C6",x"C4",x"53",x"E2",x"C2",x"F7",x"7A", -- 0x1428
		x"CE",x"74",x"04",x"A9",x"7E",x"84",x"1E",x"4F", -- 0x1430
		x"24",x"8E",x"1B",x"9E",x"7A",x"85",x"D9",x"94", -- 0x1438
		x"DB",x"CD",x"F8",x"74",x"04",x"C2",x"35",x"E1", -- 0x1440
		x"89",x"7A",x"B4",x"6C",x"3D",x"AD",x"67",x"0D", -- 0x1448
		x"A1",x"6B",x"36",x"9F",x"6F",x"54",x"EE",x"93", -- 0x1450
		x"62",x"89",x"B2",x"DC",x"0F",x"8C",x"F0",x"6A", -- 0x1458
		x"D9",x"69",x"5F",x"5E",x"2D",x"14",x"BF",x"36", -- 0x1460
		x"8E",x"74",x"23",x"CC",x"A1",x"8A",x"59",x"43", -- 0x1468
		x"75",x"8F",x"E3",x"E4",x"63",x"52",x"F7",x"C5", -- 0x1470
		x"DC",x"AA",x"22",x"6B",x"B6",x"92",x"D6",x"11", -- 0x1478
		x"FC",x"B5",x"6F",x"A9",x"C9",x"2F",x"DF",x"59", -- 0x1480
		x"A3",x"03",x"26",x"C5",x"0D",x"7F",x"09",x"82", -- 0x1488
		x"8E",x"6C",x"67",x"F1",x"BF",x"DF",x"37",x"9C", -- 0x1490
		x"0A",x"59",x"08",x"C1",x"EB",x"5E",x"D2",x"68", -- 0x1498
		x"14",x"42",x"12",x"DE",x"F0",x"F2",x"B7",x"14", -- 0x14A0
		x"75",x"DD",x"D9",x"83",x"DC",x"E3",x"06",x"6B", -- 0x14A8
		x"50",x"6E",x"DC",x"10",x"4E",x"14",x"2C",x"D7", -- 0x14B0
		x"EC",x"35",x"99",x"58",x"13",x"EB",x"C1",x"A7", -- 0x14B8
		x"2E",x"D3",x"06",x"9E",x"46",x"BD",x"B3",x"BC", -- 0x14C0
		x"1B",x"8D",x"40",x"77",x"F0",x"46",x"E2",x"C1", -- 0x14C8
		x"34",x"3F",x"51",x"02",x"53",x"7E",x"DA",x"BF", -- 0x14D0
		x"33",x"74",x"18",x"46",x"61",x"D9",x"6D",x"0F", -- 0x14D8
		x"2E",x"73",x"2E",x"74",x"31",x"E1",x"31",x"CB", -- 0x14E0
		x"EE",x"71",x"43",x"60",x"B8",x"A5",x"22",x"EC", -- 0x14E8
		x"E4",x"73",x"6F",x"B7",x"F1",x"4A",x"77",x"A4", -- 0x14F0
		x"3E",x"90",x"6B",x"1F",x"6A",x"D8",x"AE",x"98", -- 0x14F8
		x"4D",x"DC",x"8D",x"FD",x"3E",x"BE",x"CA",x"2D", -- 0x1500
		x"31",x"0E",x"8D",x"69",x"34",x"2F",x"D5",x"19", -- 0x1508
		x"A3",x"45",x"D1",x"15",x"8F",x"49",x"BA",x"4E", -- 0x1510
		x"D9",x"26",x"6D",x"C4",x"FE",x"1C",x"DC",x"CB", -- 0x1518
		x"F8",x"6A",x"4A",x"37",x"A9",x"15",x"E4",x"DA", -- 0x1520
		x"A2",x"72",x"C3",x"D6",x"22",x"99",x"70",x"C5", -- 0x1528
		x"5F",x"42",x"DA",x"6E",x"0B",x"15",x"BC",x"65", -- 0x1530
		x"3B",x"2B",x"2A",x"BA",x"47",x"86",x"06",x"C0", -- 0x1538
		x"71",x"50",x"F7",x"1B",x"65",x"DC",x"75",x"88", -- 0x1540
		x"CF",x"39",x"DE",x"F1",x"52",x"4F",x"37",x"31", -- 0x1548
		x"11",x"12",x"A0",x"1D",x"28",x"DC",x"02",x"E2", -- 0x1550
		x"87",x"AB",x"1D",x"CF",x"32",x"24",x"90",x"23", -- 0x1558
		x"74",x"08",x"3E",x"5A",x"65",x"B3",x"62",x"B4", -- 0x1560
		x"6C",x"41",x"26",x"3F",x"11",x"5D",x"EF",x"22", -- 0x1568
		x"EE",x"10",x"BE",x"96",x"ED",x"C0",x"F9",x"75", -- 0x1570
		x"6C",x"17",x"C4",x"1F",x"BA",x"D4",x"42",x"30", -- 0x1578
		x"DD",x"81",x"0A",x"C2",x"B4",x"EB",x"77",x"A1", -- 0x1580
		x"2D",x"9D",x"E0",x"3E",x"7A",x"D0",x"E0",x"69", -- 0x1588
		x"E1",x"9F",x"80",x"4F",x"E0",x"7A",x"44",x"4D", -- 0x1590
		x"91",x"0A",x"EB",x"CC",x"DE",x"2F",x"7C",x"3C", -- 0x1598
		x"30",x"86",x"7E",x"E4",x"72",x"75",x"86",x"1F", -- 0x15A0
		x"13",x"E6",x"DD",x"0D",x"38",x"BE",x"F6",x"99", -- 0x15A8
		x"DD",x"77",x"68",x"BE",x"F1",x"AC",x"8C",x"03", -- 0x15B0
		x"B6",x"78",x"CF",x"16",x"27",x"4C",x"D1",x"57", -- 0x15B8
		x"52",x"D0",x"BC",x"44",x"46",x"C2",x"64",x"D9", -- 0x15C0
		x"AA",x"C1",x"E6",x"62",x"00",x"DD",x"7B",x"DD", -- 0x15C8
		x"D4",x"E3",x"1D",x"C6",x"10",x"29",x"4A",x"47", -- 0x15D0
		x"21",x"99",x"DC",x"49",x"66",x"AE",x"20",x"B8", -- 0x15D8
		x"FE",x"DC",x"FD",x"46",x"A0",x"E1",x"20",x"CA", -- 0x15E0
		x"23",x"86",x"AC",x"23",x"65",x"28",x"01",x"3A", -- 0x15E8
		x"8B",x"9D",x"81",x"9B",x"C6",x"4B",x"E2",x"68", -- 0x15F0
		x"E4",x"3F",x"B1",x"4B",x"EE",x"D1",x"84",x"6D", -- 0x15F8
		x"2F",x"02",x"B3",x"CF",x"E3",x"53",x"9A",x"86", -- 0x1600
		x"DA",x"C6",x"A9",x"40",x"EE",x"2A",x"F9",x"F9", -- 0x1608
		x"C8",x"FA",x"15",x"0F",x"46",x"78",x"77",x"AB", -- 0x1610
		x"B7",x"A8",x"F6",x"26",x"FA",x"FA",x"94",x"2A", -- 0x1618
		x"FC",x"48",x"F9",x"E0",x"9C",x"14",x"E6",x"F6", -- 0x1620
		x"DA",x"90",x"37",x"49",x"BB",x"B0",x"43",x"84", -- 0x1628
		x"AC",x"D7",x"13",x"72",x"50",x"8B",x"1E",x"09", -- 0x1630
		x"34",x"95",x"2F",x"2F",x"90",x"43",x"59",x"8E", -- 0x1638
		x"0C",x"D2",x"EE",x"A8",x"66",x"D6",x"1F",x"C0", -- 0x1640
		x"E6",x"56",x"0A",x"A2",x"86",x"CC",x"A6",x"B2", -- 0x1648
		x"25",x"BA",x"26",x"75",x"46",x"C3",x"FD",x"F9", -- 0x1650
		x"D8",x"2E",x"2A",x"E9",x"F0",x"03",x"78",x"FC", -- 0x1658
		x"56",x"E6",x"25",x"3C",x"3D",x"44",x"FD",x"25", -- 0x1660
		x"1A",x"87",x"47",x"A1",x"D4",x"EE",x"54",x"F9", -- 0x1668
		x"A9",x"F9",x"6F",x"6F",x"3E",x"6E",x"69",x"96", -- 0x1670
		x"1C",x"13",x"80",x"0D",x"96",x"78",x"8A",x"EC", -- 0x1678
		x"DF",x"AF",x"29",x"1D",x"F4",x"A6",x"C1",x"0F", -- 0x1680
		x"2F",x"0A",x"30",x"83",x"F8",x"05",x"7D",x"A2", -- 0x1688
		x"7E",x"6C",x"91",x"BC",x"5A",x"FA",x"D3",x"F5", -- 0x1690
		x"0F",x"54",x"04",x"A5",x"CD",x"0E",x"12",x"AD", -- 0x1698
		x"BD",x"BA",x"4A",x"32",x"62",x"0D",x"42",x"11", -- 0x16A0
		x"96",x"F1",x"94",x"8F",x"F6",x"91",x"B1",x"76", -- 0x16A8
		x"FD",x"43",x"B2",x"D8",x"3E",x"86",x"CE",x"CC", -- 0x16B0
		x"DB",x"52",x"72",x"29",x"60",x"04",x"56",x"1F", -- 0x16B8
		x"BF",x"20",x"51",x"A1",x"AC",x"13",x"B2",x"43", -- 0x16C0
		x"06",x"C6",x"D2",x"7C",x"58",x"04",x"F2",x"D5", -- 0x16C8
		x"C6",x"26",x"AE",x"85",x"AC",x"7E",x"52",x"08", -- 0x16D0
		x"50",x"45",x"B0",x"B1",x"49",x"07",x"50",x"88", -- 0x16D8
		x"A7",x"A1",x"2A",x"54",x"35",x"DC",x"98",x"BA", -- 0x16E0
		x"23",x"EA",x"37",x"FA",x"EF",x"AA",x"51",x"B6", -- 0x16E8
		x"D0",x"00",x"3C",x"FC",x"FD",x"0F",x"06",x"4F", -- 0x16F0
		x"54",x"36",x"80",x"1D",x"BD",x"D0",x"A6",x"65", -- 0x16F8
		x"F1",x"D0",x"B9",x"27",x"2E",x"52",x"61",x"D0", -- 0x1700
		x"BD",x"99",x"CC",x"2D",x"C3",x"1E",x"E3",x"94", -- 0x1708
		x"9D",x"A0",x"11",x"1C",x"2F",x"96",x"6B",x"03", -- 0x1710
		x"CD",x"6B",x"20",x"8B",x"3C",x"46",x"F0",x"2E", -- 0x1718
		x"97",x"2A",x"D5",x"45",x"FC",x"37",x"16",x"BA", -- 0x1720
		x"D0",x"62",x"E7",x"14",x"80",x"4B",x"28",x"1F", -- 0x1728
		x"6B",x"3A",x"BA",x"9A",x"D0",x"26",x"9D",x"1E", -- 0x1730
		x"11",x"3E",x"A9",x"4D",x"04",x"1A",x"7B",x"9B", -- 0x1738
		x"45",x"51",x"E0",x"42",x"89",x"77",x"FC",x"D9", -- 0x1740
		x"D9",x"64",x"6E",x"5B",x"AF",x"96",x"F9",x"1C", -- 0x1748
		x"D0",x"B4",x"B6",x"22",x"5A",x"D4",x"40",x"6B", -- 0x1750
		x"92",x"6A",x"38",x"96",x"84",x"33",x"33",x"49", -- 0x1758
		x"85",x"93",x"8B",x"8E",x"0B",x"08",x"E7",x"65", -- 0x1760
		x"6C",x"56",x"C0",x"9C",x"6D",x"3A",x"B8",x"BD", -- 0x1768
		x"6E",x"EE",x"DF",x"48",x"C3",x"A0",x"33",x"56", -- 0x1770
		x"8A",x"6B",x"6D",x"8E",x"1E",x"A0",x"D8",x"A3", -- 0x1778
		x"B3",x"E3",x"B1",x"3F",x"6C",x"1A",x"A4",x"58", -- 0x1780
		x"EF",x"65",x"F4",x"5D",x"1F",x"AD",x"1C",x"0D", -- 0x1788
		x"9D",x"7B",x"D4",x"E0",x"9B",x"08",x"B7",x"26", -- 0x1790
		x"F2",x"25",x"B5",x"11",x"45",x"0E",x"35",x"F8", -- 0x1798
		x"71",x"66",x"38",x"DD",x"80",x"DC",x"37",x"71", -- 0x17A0
		x"C1",x"2C",x"CE",x"60",x"DA",x"6A",x"EC",x"F7", -- 0x17A8
		x"E6",x"C1",x"58",x"82",x"C9",x"10",x"29",x"3C", -- 0x17B0
		x"B4",x"5E",x"CD",x"79",x"6C",x"03",x"73",x"5D", -- 0x17B8
		x"E8",x"2B",x"3C",x"6A",x"88",x"F2",x"5B",x"C9", -- 0x17C0
		x"1F",x"A9",x"AA",x"79",x"15",x"97",x"F0",x"7B", -- 0x17C8
		x"5A",x"4A",x"7D",x"A3",x"D9",x"A6",x"60",x"0F", -- 0x17D0
		x"05",x"2E",x"88",x"F0",x"B0",x"7B",x"4F",x"99", -- 0x17D8
		x"27",x"0B",x"83",x"AF",x"FD",x"DE",x"F8",x"9C", -- 0x17E0
		x"89",x"23",x"96",x"1E",x"BB",x"87",x"99",x"95", -- 0x17E8
		x"51",x"96",x"B8",x"AB",x"3E",x"19",x"BA",x"C2", -- 0x17F0
		x"C6",x"43",x"34",x"F6",x"BF",x"03",x"91",x"E6", -- 0x17F8
		x"0E",x"15",x"16",x"8B",x"74",x"0F",x"A7",x"FD", -- 0x1800
		x"33",x"3E",x"9B",x"6E",x"46",x"35",x"83",x"97", -- 0x1808
		x"CB",x"3C",x"C2",x"89",x"D5",x"7D",x"CC",x"1C", -- 0x1810
		x"C1",x"01",x"14",x"81",x"04",x"A5",x"E7",x"91", -- 0x1818
		x"3A",x"FD",x"9C",x"AE",x"8C",x"44",x"2C",x"3F", -- 0x1820
		x"03",x"C7",x"AD",x"49",x"FC",x"31",x"60",x"49", -- 0x1828
		x"ED",x"24",x"52",x"43",x"A1",x"1F",x"5F",x"63", -- 0x1830
		x"9F",x"73",x"64",x"23",x"98",x"4C",x"B4",x"D3", -- 0x1838
		x"C9",x"D0",x"02",x"57",x"16",x"2F",x"96",x"19", -- 0x1840
		x"F6",x"45",x"E1",x"74",x"F5",x"42",x"BD",x"63", -- 0x1848
		x"66",x"8F",x"A6",x"88",x"AF",x"07",x"6B",x"CE", -- 0x1850
		x"F9",x"D0",x"F2",x"93",x"9C",x"A7",x"E6",x"67", -- 0x1858
		x"79",x"E8",x"BE",x"0F",x"18",x"55",x"A7",x"10", -- 0x1860
		x"1A",x"89",x"84",x"90",x"CB",x"C1",x"F3",x"B2", -- 0x1868
		x"D0",x"1B",x"3B",x"00",x"A1",x"A6",x"CF",x"9B", -- 0x1870
		x"F6",x"C2",x"AE",x"14",x"E9",x"15",x"7B",x"E2", -- 0x1878
		x"FE",x"B9",x"F1",x"96",x"0F",x"19",x"A6",x"A9", -- 0x1880
		x"A2",x"AA",x"B9",x"6F",x"EB",x"2D",x"A1",x"3D", -- 0x1888
		x"48",x"5C",x"3D",x"69",x"82",x"0D",x"85",x"7A", -- 0x1890
		x"4F",x"34",x"0E",x"B9",x"4A",x"89",x"9C",x"C8", -- 0x1898
		x"43",x"0F",x"5F",x"D1",x"28",x"86",x"FA",x"CB", -- 0x18A0
		x"B0",x"B4",x"BA",x"1D",x"E2",x"DB",x"5A",x"AA", -- 0x18A8
		x"38",x"97",x"94",x"BA",x"25",x"1A",x"B4",x"F3", -- 0x18B0
		x"CD",x"C2",x"AD",x"97",x"CB",x"4B",x"60",x"8E", -- 0x18B8
		x"D9",x"40",x"61",x"02",x"C6",x"DB",x"4D",x"F6", -- 0x18C0
		x"91",x"87",x"14",x"F3",x"63",x"6E",x"1E",x"1B", -- 0x18C8
		x"86",x"B2",x"56",x"AB",x"4C",x"8A",x"9F",x"1B", -- 0x18D0
		x"CD",x"4E",x"B2",x"99",x"19",x"93",x"29",x"F2", -- 0x18D8
		x"53",x"0A",x"74",x"99",x"E5",x"C2",x"90",x"F6", -- 0x18E0
		x"C9",x"A5",x"6A",x"2E",x"93",x"89",x"C8",x"1A", -- 0x18E8
		x"BB",x"1F",x"45",x"09",x"AA",x"E5",x"A3",x"78", -- 0x18F0
		x"B3",x"D5",x"91",x"CC",x"E8",x"3A",x"3F",x"3C", -- 0x18F8
		x"44",x"B3",x"D5",x"AA",x"F5",x"67",x"21",x"C0", -- 0x1900
		x"8C",x"8C",x"EE",x"20",x"95",x"37",x"BA",x"D0", -- 0x1908
		x"57",x"00",x"D9",x"02",x"65",x"FC",x"F9",x"19", -- 0x1910
		x"D3",x"8B",x"65",x"BC",x"C6",x"A4",x"F9",x"8A", -- 0x1918
		x"D8",x"4F",x"35",x"CE",x"36",x"57",x"8F",x"C2", -- 0x1920
		x"63",x"FD",x"63",x"78",x"36",x"1E",x"49",x"0D", -- 0x1928
		x"9D",x"24",x"0F",x"04",x"A0",x"88",x"1D",x"74", -- 0x1930
		x"14",x"03",x"B1",x"DA",x"27",x"AB",x"E5",x"00", -- 0x1938
		x"7A",x"1B",x"4F",x"B1",x"F1",x"5E",x"74",x"D4", -- 0x1940
		x"5D",x"57",x"4D",x"13",x"F4",x"97",x"20",x"93", -- 0x1948
		x"3B",x"AE",x"97",x"DB",x"37",x"34",x"D0",x"4B", -- 0x1950
		x"B6",x"82",x"A6",x"DE",x"AD",x"8C",x"5E",x"28", -- 0x1958
		x"27",x"AD",x"D9",x"99",x"0D",x"CE",x"6E",x"E9", -- 0x1960
		x"26",x"BC",x"FC",x"1C",x"D3",x"9C",x"2F",x"0F", -- 0x1968
		x"4B",x"46",x"6A",x"82",x"F9",x"3B",x"4D",x"B1", -- 0x1970
		x"BD",x"73",x"10",x"6B",x"7F",x"6E",x"14",x"A7", -- 0x1978
		x"9C",x"ED",x"41",x"A9",x"BC",x"2F",x"13",x"E3", -- 0x1980
		x"6B",x"8F",x"7F",x"3F",x"2C",x"2E",x"CD",x"F6", -- 0x1988
		x"74",x"39",x"F8",x"ED",x"F3",x"C5",x"9F",x"32", -- 0x1990
		x"3A",x"AF",x"1D",x"B9",x"9E",x"31",x"E0",x"3B", -- 0x1998
		x"20",x"A1",x"64",x"5C",x"D1",x"77",x"BF",x"BC", -- 0x19A0
		x"86",x"3F",x"FC",x"32",x"EC",x"4A",x"29",x"E0", -- 0x19A8
		x"03",x"A1",x"CF",x"F7",x"67",x"EE",x"A9",x"21", -- 0x19B0
		x"9F",x"C6",x"DB",x"BD",x"F8",x"3C",x"F8",x"98", -- 0x19B8
		x"DE",x"5D",x"F4",x"B0",x"54",x"B5",x"EC",x"DA", -- 0x19C0
		x"74",x"E9",x"0D",x"E1",x"B4",x"B5",x"C2",x"B7", -- 0x19C8
		x"57",x"12",x"2F",x"BE",x"02",x"D8",x"E0",x"21", -- 0x19D0
		x"A0",x"3C",x"DE",x"19",x"78",x"D7",x"31",x"D6", -- 0x19D8
		x"B4",x"26",x"07",x"09",x"5B",x"F4",x"E3",x"50", -- 0x19E0
		x"DE",x"70",x"32",x"13",x"26",x"74",x"CB",x"7D", -- 0x19E8
		x"87",x"FA",x"BB",x"89",x"D4",x"1C",x"AA",x"F4", -- 0x19F0
		x"D7",x"89",x"0E",x"D0",x"61",x"BE",x"A7",x"16", -- 0x19F8
		x"64",x"AF",x"9E",x"C0",x"A4",x"02",x"90",x"03", -- 0x1A00
		x"72",x"42",x"17",x"98",x"B6",x"62",x"95",x"3E", -- 0x1A08
		x"5D",x"51",x"C7",x"B1",x"ED",x"72",x"A6",x"C5", -- 0x1A10
		x"7B",x"34",x"96",x"5C",x"F2",x"3F",x"F1",x"D7", -- 0x1A18
		x"6E",x"90",x"18",x"13",x"92",x"A8",x"95",x"05", -- 0x1A20
		x"EA",x"AC",x"1D",x"A1",x"8E",x"B2",x"60",x"EC", -- 0x1A28
		x"84",x"28",x"1E",x"F1",x"1B",x"C5",x"B7",x"16", -- 0x1A30
		x"79",x"4F",x"73",x"EC",x"0E",x"65",x"C4",x"7C", -- 0x1A38
		x"76",x"DC",x"0F",x"88",x"05",x"A4",x"0E",x"EF", -- 0x1A40
		x"D1",x"2B",x"11",x"60",x"5E",x"F0",x"4D",x"62", -- 0x1A48
		x"99",x"6C",x"54",x"34",x"B1",x"0C",x"4A",x"AA", -- 0x1A50
		x"DA",x"BD",x"97",x"E8",x"A3",x"5C",x"E4",x"99", -- 0x1A58
		x"B8",x"F3",x"22",x"BD",x"99",x"30",x"2D",x"6B", -- 0x1A60
		x"DB",x"BE",x"4B",x"3A",x"AF",x"19",x"1C",x"49", -- 0x1A68
		x"05",x"70",x"7D",x"B6",x"FB",x"48",x"61",x"57", -- 0x1A70
		x"85",x"F9",x"BF",x"29",x"D5",x"A5",x"42",x"0F", -- 0x1A78
		x"19",x"65",x"CC",x"B2",x"15",x"7A",x"9D",x"F0", -- 0x1A80
		x"39",x"E9",x"AA",x"68",x"82",x"46",x"B2",x"87", -- 0x1A88
		x"B6",x"AF",x"3E",x"33",x"F7",x"1F",x"8A",x"7E", -- 0x1A90
		x"98",x"4A",x"27",x"6F",x"6F",x"6A",x"FD",x"89", -- 0x1A98
		x"4F",x"CA",x"3C",x"E3",x"45",x"5A",x"D5",x"FD", -- 0x1AA0
		x"C3",x"00",x"67",x"46",x"47",x"99",x"CD",x"7D", -- 0x1AA8
		x"49",x"8B",x"B0",x"42",x"AA",x"BA",x"40",x"44", -- 0x1AB0
		x"06",x"67",x"33",x"75",x"51",x"31",x"7E",x"20", -- 0x1AB8
		x"7B",x"BB",x"05",x"41",x"95",x"DA",x"3F",x"D8", -- 0x1AC0
		x"5A",x"A6",x"1F",x"A1",x"40",x"6C",x"9F",x"0A", -- 0x1AC8
		x"F7",x"50",x"CB",x"22",x"8B",x"0C",x"E5",x"91", -- 0x1AD0
		x"F2",x"98",x"86",x"C4",x"49",x"06",x"E4",x"C5", -- 0x1AD8
		x"41",x"E9",x"86",x"56",x"C4",x"C5",x"2F",x"9F", -- 0x1AE0
		x"EC",x"CD",x"C0",x"AC",x"B9",x"60",x"B6",x"31", -- 0x1AE8
		x"31",x"82",x"53",x"BC",x"0E",x"B9",x"CD",x"02", -- 0x1AF0
		x"52",x"D3",x"C6",x"1C",x"59",x"AB",x"61",x"1A", -- 0x1AF8
		x"16",x"E7",x"70",x"5A",x"2D",x"1F",x"F9",x"1A", -- 0x1B00
		x"6C",x"BB",x"C7",x"26",x"1C",x"FD",x"57",x"CC", -- 0x1B08
		x"01",x"2B",x"89",x"0F",x"64",x"D6",x"90",x"B6", -- 0x1B10
		x"AB",x"D6",x"52",x"05",x"03",x"B3",x"9F",x"19", -- 0x1B18
		x"9B",x"10",x"73",x"C9",x"AF",x"6E",x"63",x"1C", -- 0x1B20
		x"A9",x"AA",x"43",x"45",x"A9",x"1A",x"13",x"2A", -- 0x1B28
		x"45",x"1C",x"39",x"A9",x"F3",x"4A",x"E0",x"9F", -- 0x1B30
		x"A0",x"33",x"24",x"A3",x"67",x"C3",x"3C",x"03", -- 0x1B38
		x"54",x"30",x"4C",x"04",x"1E",x"30",x"20",x"C7", -- 0x1B40
		x"DA",x"E2",x"0D",x"04",x"FD",x"9F",x"2E",x"C2", -- 0x1B48
		x"BC",x"E7",x"EC",x"B0",x"B1",x"CD",x"CF",x"52", -- 0x1B50
		x"80",x"73",x"76",x"E7",x"B7",x"B2",x"6B",x"0C", -- 0x1B58
		x"62",x"37",x"8F",x"80",x"67",x"AF",x"48",x"C2", -- 0x1B60
		x"93",x"D5",x"46",x"11",x"75",x"75",x"D3",x"32", -- 0x1B68
		x"DC",x"C0",x"62",x"8E",x"0E",x"32",x"60",x"0F", -- 0x1B70
		x"26",x"D6",x"76",x"DD",x"0A",x"61",x"E9",x"6C", -- 0x1B78
		x"99",x"79",x"ED",x"80",x"A8",x"B5",x"C2",x"BB", -- 0x1B80
		x"0B",x"0A",x"CC",x"81",x"FE",x"21",x"33",x"DB", -- 0x1B88
		x"61",x"16",x"E9",x"70",x"C7",x"4A",x"7F",x"ED", -- 0x1B90
		x"22",x"75",x"CB",x"2C",x"D7",x"B5",x"98",x"71", -- 0x1B98
		x"AE",x"06",x"71",x"D7",x"BC",x"35",x"93",x"C7", -- 0x1BA0
		x"BE",x"E0",x"C8",x"BD",x"81",x"7C",x"19",x"E2", -- 0x1BA8
		x"92",x"03",x"D2",x"5A",x"CC",x"D1",x"C8",x"6E", -- 0x1BB0
		x"48",x"94",x"9A",x"20",x"CA",x"B3",x"11",x"F8", -- 0x1BB8
		x"B9",x"82",x"D0",x"F5",x"37",x"E4",x"3E",x"75", -- 0x1BC0
		x"C5",x"07",x"33",x"47",x"03",x"CB",x"A9",x"95", -- 0x1BC8
		x"4E",x"7D",x"70",x"9B",x"4F",x"39",x"0A",x"97", -- 0x1BD0
		x"4D",x"25",x"B7",x"18",x"D8",x"48",x"12",x"12", -- 0x1BD8
		x"4B",x"E2",x"88",x"02",x"47",x"C6",x"78",x"0D", -- 0x1BE0
		x"4D",x"2B",x"D3",x"51",x"77",x"7E",x"66",x"C5", -- 0x1BE8
		x"7B",x"56",x"61",x"CA",x"8F",x"6C",x"E2",x"5D", -- 0x1BF0
		x"91",x"1A",x"75",x"E9",x"63",x"07",x"7B",x"AE", -- 0x1BF8
		x"EA",x"04",x"30",x"32",x"CA",x"A8",x"BF",x"19", -- 0x1C00
		x"54",x"13",x"E9",x"CB",x"11",x"50",x"91",x"8C", -- 0x1C08
		x"A7",x"73",x"D7",x"B6",x"5F",x"BA",x"14",x"F0", -- 0x1C10
		x"D4",x"8A",x"5A",x"B7",x"11",x"D5",x"E5",x"FB", -- 0x1C18
		x"5A",x"17",x"AE",x"A4",x"BF",x"ED",x"3D",x"14", -- 0x1C20
		x"80",x"27",x"DF",x"92",x"78",x"F1",x"9E",x"20", -- 0x1C28
		x"65",x"76",x"56",x"44",x"B0",x"6B",x"B4",x"86", -- 0x1C30
		x"75",x"0F",x"BD",x"86",x"64",x"A4",x"03",x"3E", -- 0x1C38
		x"BB",x"31",x"E3",x"7B",x"9E",x"21",x"10",x"1F", -- 0x1C40
		x"49",x"6F",x"31",x"C1",x"E0",x"D0",x"61",x"C5", -- 0x1C48
		x"C6",x"B7",x"0A",x"78",x"A2",x"BE",x"7E",x"18", -- 0x1C50
		x"CD",x"BB",x"1F",x"B2",x"60",x"22",x"F0",x"1C", -- 0x1C58
		x"D2",x"54",x"18",x"71",x"76",x"A7",x"90",x"BF", -- 0x1C60
		x"17",x"C2",x"01",x"F8",x"13",x"E1",x"3E",x"59", -- 0x1C68
		x"99",x"49",x"51",x"3D",x"08",x"CF",x"D4",x"56", -- 0x1C70
		x"8C",x"F3",x"88",x"6C",x"95",x"79",x"89",x"68", -- 0x1C78
		x"4E",x"A1",x"D9",x"C4",x"49",x"EA",x"04",x"DF", -- 0x1C80
		x"AD",x"84",x"58",x"40",x"66",x"97",x"99",x"7F", -- 0x1C88
		x"E0",x"EB",x"3C",x"68",x"3B",x"12",x"BE",x"47", -- 0x1C90
		x"85",x"C6",x"B4",x"1C",x"C0",x"BD",x"84",x"0F", -- 0x1C98
		x"DE",x"5F",x"D3",x"A7",x"4A",x"D7",x"87",x"77", -- 0x1CA0
		x"5C",x"60",x"37",x"42",x"F7",x"D0",x"C1",x"58", -- 0x1CA8
		x"3C",x"FE",x"C0",x"78",x"90",x"00",x"3F",x"16", -- 0x1CB0
		x"C6",x"F3",x"32",x"87",x"31",x"37",x"96",x"10", -- 0x1CB8
		x"16",x"6A",x"B7",x"DF",x"C1",x"BF",x"D6",x"9D", -- 0x1CC0
		x"20",x"0E",x"5F",x"18",x"5E",x"22",x"70",x"9B", -- 0x1CC8
		x"A0",x"B0",x"93",x"31",x"B0",x"D2",x"47",x"F7", -- 0x1CD0
		x"47",x"F9",x"7F",x"78",x"31",x"96",x"89",x"C6", -- 0x1CD8
		x"80",x"41",x"A6",x"43",x"80",x"7D",x"60",x"A0", -- 0x1CE0
		x"0B",x"C0",x"B8",x"69",x"62",x"A8",x"05",x"03", -- 0x1CE8
		x"D9",x"98",x"34",x"0A",x"EB",x"FA",x"02",x"33", -- 0x1CF0
		x"F4",x"82",x"AB",x"A5",x"98",x"B4",x"EB",x"19", -- 0x1CF8
		x"76",x"92",x"DB",x"F6",x"8F",x"3D",x"98",x"1A", -- 0x1D00
		x"7D",x"D0",x"84",x"DF",x"F9",x"09",x"E2",x"D3", -- 0x1D08
		x"A2",x"96",x"DD",x"8E",x"91",x"E0",x"41",x"07", -- 0x1D10
		x"E2",x"EC",x"2C",x"7B",x"22",x"19",x"94",x"98", -- 0x1D18
		x"2B",x"F0",x"8F",x"3B",x"2E",x"28",x"55",x"2B", -- 0x1D20
		x"79",x"59",x"0B",x"73",x"63",x"6D",x"47",x"85", -- 0x1D28
		x"83",x"A4",x"14",x"15",x"85",x"D4",x"9B",x"E7", -- 0x1D30
		x"C1",x"C8",x"E2",x"E3",x"61",x"F7",x"FB",x"0C", -- 0x1D38
		x"E8",x"8C",x"47",x"17",x"34",x"1D",x"C1",x"AD", -- 0x1D40
		x"76",x"CC",x"A0",x"59",x"B9",x"E7",x"DE",x"3D", -- 0x1D48
		x"8D",x"F2",x"D1",x"92",x"C7",x"6E",x"FA",x"0A", -- 0x1D50
		x"B6",x"DD",x"6D",x"97",x"D5",x"6A",x"A3",x"BE", -- 0x1D58
		x"76",x"6B",x"55",x"2A",x"08",x"17",x"58",x"FD", -- 0x1D60
		x"63",x"F8",x"58",x"9C",x"61",x"37",x"59",x"6E", -- 0x1D68
		x"AA",x"2C",x"01",x"F1",x"1A",x"FB",x"FB",x"50", -- 0x1D70
		x"5A",x"E9",x"E7",x"30",x"D3",x"0B",x"6F",x"4A", -- 0x1D78
		x"76",x"C4",x"74",x"FD",x"5C",x"4C",x"FC",x"3F", -- 0x1D80
		x"46",x"55",x"DC",x"A7",x"0C",x"36",x"16",x"B6", -- 0x1D88
		x"E1",x"96",x"A9",x"FB",x"13",x"25",x"4C",x"6D", -- 0x1D90
		x"8E",x"34",x"1D",x"62",x"BF",x"8C",x"2C",x"36", -- 0x1D98
		x"52",x"21",x"B4",x"2E",x"6D",x"B1",x"6D",x"B3", -- 0x1DA0
		x"86",x"C9",x"DA",x"92",x"01",x"F0",x"C9",x"E2", -- 0x1DA8
		x"08",x"73",x"5F",x"1B",x"18",x"AB",x"08",x"A7", -- 0x1DB0
		x"60",x"25",x"0A",x"20",x"B2",x"B6",x"D5",x"84", -- 0x1DB8
		x"D7",x"0A",x"B2",x"45",x"BB",x"9F",x"79",x"C1", -- 0x1DC0
		x"6A",x"54",x"D4",x"EA",x"C5",x"1E",x"CD",x"CD", -- 0x1DC8
		x"11",x"AC",x"68",x"29",x"59",x"70",x"D0",x"39", -- 0x1DD0
		x"95",x"5B",x"D8",x"C7",x"12",x"2E",x"CB",x"69", -- 0x1DD8
		x"39",x"7E",x"2E",x"74",x"9E",x"A7",x"37",x"09", -- 0x1DE0
		x"7C",x"8B",x"F3",x"42",x"A9",x"41",x"8F",x"BA", -- 0x1DE8
		x"EE",x"F7",x"63",x"C7",x"E7",x"B4",x"80",x"FC", -- 0x1DF0
		x"10",x"59",x"C5",x"A1",x"87",x"91",x"8A",x"C0", -- 0x1DF8
		x"90",x"B8",x"36",x"2F",x"61",x"EC",x"B7",x"DD", -- 0x1E00
		x"F7",x"2B",x"9F",x"21",x"EB",x"2F",x"DB",x"DA", -- 0x1E08
		x"27",x"BE",x"22",x"0F",x"73",x"A2",x"0C",x"03", -- 0x1E10
		x"7B",x"51",x"A4",x"04",x"63",x"2F",x"44",x"F3", -- 0x1E18
		x"68",x"F9",x"A2",x"C9",x"E6",x"D9",x"27",x"5E", -- 0x1E20
		x"05",x"C6",x"7F",x"F0",x"F5",x"DA",x"4C",x"9C", -- 0x1E28
		x"9A",x"ED",x"2B",x"0E",x"11",x"B6",x"91",x"8C", -- 0x1E30
		x"09",x"36",x"10",x"EB",x"E5",x"55",x"5F",x"4E", -- 0x1E38
		x"CE",x"02",x"97",x"36",x"5B",x"BE",x"94",x"60", -- 0x1E40
		x"05",x"15",x"D0",x"7A",x"6F",x"9C",x"17",x"0A", -- 0x1E48
		x"8B",x"42",x"98",x"9C",x"78",x"2A",x"A8",x"01", -- 0x1E50
		x"DF",x"B9",x"EC",x"45",x"8E",x"4C",x"93",x"5D", -- 0x1E58
		x"CD",x"AA",x"93",x"29",x"E8",x"A8",x"09",x"ED", -- 0x1E60
		x"BD",x"DA",x"68",x"AC",x"77",x"FE",x"B7",x"82", -- 0x1E68
		x"C0",x"50",x"9E",x"3A",x"F9",x"48",x"3B",x"D9", -- 0x1E70
		x"81",x"29",x"20",x"10",x"F4",x"33",x"EC",x"C3", -- 0x1E78
		x"5E",x"01",x"EC",x"47",x"A9",x"F6",x"B5",x"E6", -- 0x1E80
		x"51",x"9D",x"93",x"48",x"9D",x"4B",x"CB",x"5E", -- 0x1E88
		x"1B",x"E9",x"98",x"94",x"32",x"D4",x"6F",x"B3", -- 0x1E90
		x"7D",x"0F",x"43",x"72",x"42",x"31",x"36",x"20", -- 0x1E98
		x"32",x"A3",x"68",x"5B",x"9A",x"1E",x"42",x"6B", -- 0x1EA0
		x"BB",x"D5",x"B3",x"D8",x"A1",x"FE",x"38",x"3C", -- 0x1EA8
		x"E9",x"D0",x"D1",x"9B",x"25",x"C0",x"CF",x"A2", -- 0x1EB0
		x"CF",x"13",x"16",x"91",x"C3",x"CB",x"B2",x"75", -- 0x1EB8
		x"6F",x"9A",x"D0",x"89",x"38",x"13",x"F4",x"F3", -- 0x1EC0
		x"69",x"29",x"4D",x"8A",x"28",x"85",x"C6",x"91", -- 0x1EC8
		x"D5",x"18",x"AD",x"FB",x"D8",x"7D",x"1E",x"28", -- 0x1ED0
		x"10",x"B3",x"BA",x"D4",x"80",x"EC",x"4A",x"6F", -- 0x1ED8
		x"87",x"1C",x"F9",x"BF",x"AE",x"EE",x"33",x"18", -- 0x1EE0
		x"18",x"80",x"A2",x"C0",x"85",x"E9",x"D1",x"5C", -- 0x1EE8
		x"02",x"7F",x"58",x"5B",x"FC",x"76",x"83",x"0E", -- 0x1EF0
		x"AA",x"BD",x"62",x"2B",x"2A",x"AC",x"9A",x"B1", -- 0x1EF8
		x"48",x"14",x"F0",x"F7",x"04",x"A4",x"8F",x"9B", -- 0x1F00
		x"25",x"33",x"DB",x"AB",x"9C",x"AE",x"08",x"9E", -- 0x1F08
		x"2E",x"DF",x"F9",x"AB",x"D5",x"FD",x"39",x"80", -- 0x1F10
		x"3B",x"9B",x"2B",x"66",x"C7",x"46",x"18",x"90", -- 0x1F18
		x"5A",x"89",x"08",x"DD",x"2E",x"97",x"7A",x"D2", -- 0x1F20
		x"4A",x"D5",x"7E",x"E6",x"84",x"06",x"86",x"33", -- 0x1F28
		x"65",x"00",x"DE",x"BB",x"7D",x"97",x"3C",x"B9", -- 0x1F30
		x"33",x"E7",x"20",x"7A",x"2E",x"B7",x"0B",x"88", -- 0x1F38
		x"41",x"92",x"67",x"EE",x"2B",x"61",x"C2",x"75", -- 0x1F40
		x"37",x"C0",x"5D",x"3C",x"47",x"63",x"6F",x"AC", -- 0x1F48
		x"E2",x"CD",x"68",x"61",x"65",x"25",x"1B",x"98", -- 0x1F50
		x"0D",x"3B",x"92",x"BA",x"72",x"1E",x"C2",x"B4", -- 0x1F58
		x"B0",x"A9",x"23",x"DB",x"0B",x"E5",x"D1",x"C2", -- 0x1F60
		x"A7",x"AE",x"FE",x"EE",x"91",x"6E",x"1B",x"74", -- 0x1F68
		x"3C",x"04",x"55",x"21",x"29",x"EF",x"B9",x"B5", -- 0x1F70
		x"2B",x"CB",x"70",x"1E",x"E9",x"B2",x"52",x"1B", -- 0x1F78
		x"5D",x"75",x"76",x"E7",x"5C",x"48",x"AA",x"83", -- 0x1F80
		x"76",x"29",x"F1",x"87",x"17",x"0D",x"7C",x"D2", -- 0x1F88
		x"11",x"D1",x"F3",x"B9",x"C2",x"2D",x"6F",x"6D", -- 0x1F90
		x"F9",x"5F",x"8B",x"63",x"13",x"DD",x"7E",x"EF", -- 0x1F98
		x"D3",x"F5",x"D7",x"30",x"BD",x"03",x"33",x"B4", -- 0x1FA0
		x"2C",x"25",x"3C",x"44",x"B1",x"B8",x"17",x"43", -- 0x1FA8
		x"0B",x"8B",x"FC",x"CD",x"B8",x"EC",x"BA",x"B2", -- 0x1FB0
		x"4C",x"47",x"17",x"DE",x"A4",x"15",x"CE",x"78", -- 0x1FB8
		x"8A",x"27",x"28",x"49",x"2A",x"DA",x"7D",x"56", -- 0x1FC0
		x"00",x"B9",x"1A",x"32",x"F2",x"B1",x"75",x"FD", -- 0x1FC8
		x"3D",x"F1",x"4B",x"F5",x"DE",x"06",x"29",x"2C", -- 0x1FD0
		x"CC",x"BF",x"8A",x"72",x"D4",x"5A",x"6A",x"60", -- 0x1FD8
		x"81",x"13",x"29",x"2B",x"ED",x"26",x"01",x"6E", -- 0x1FE0
		x"5F",x"1C",x"A0",x"52",x"4D",x"95",x"CF",x"8A", -- 0x1FE8
		x"87",x"1B",x"00",x"67",x"22",x"A8",x"93",x"6E", -- 0x1FF0
		x"68",x"9D",x"E0",x"BD",x"F7",x"CB",x"9D",x"F8"  -- 0x1FF8
	);
	attribute ram_style : string;
	attribute ram_style of ROM : signal is "block";

begin

	p_rom : process(CLK,ADDR)
	begin
		if (rising_edge(CLK)) then
			DATA <= ROM(to_integer(unsigned(ADDR)));
		 end if;
	end process;
end RTL;
