library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CartTable is
   port(clk: in std_logic;
        d: out std_logic_vector(10 downto 0);  -- rom config
        c: out std_logic_vector(6 downto 0);   -- card max
        a: in std_logic_vector(6 downto 0));   -- card control
end CartTable;

-- Bank switching(3 downto 1);
-- Superchip(0);

architecture arch of CartTable is
   type rom_type is array (0 to 127) of std_logic_vector(10 downto 0);
   signal rom: rom_type := (
      "00000000000",
      "00000010000",
      "00000100010",
      "00001000010",
      "00001100010",
      "00010000100",
      "00011000101",
      "00100000011",
      "00100100010",
      "00101000101",
      "00110000000",
      "00110010000",
      "00110100000",
      "00110110000",
      "00111000010",
      "00111100010",
      "01000001000",
      "01000101000",
      "01001000000",
      "01001010000",
      "01001100000",
      "01001110000",
      "01010000101",
      "01011000010",
      "01011100010",
      "01100000010",
      "01100100010",
      "01101000100",
      "01110000000",
      "01110010000",
      "01110100000",
      "01110110000",
      "01111000100",
      "10000000010",
      "10000100010",
      "10001000000",
      "10001010000",
      "10001100010",
      "10010000100",
      "10011000010",
      "10011100010",
      "10100000100",
      "10101000010",
      "10101100010",
      "10110000100",
      "10111001010",
      "10111101010",
      "11000001010",
      "11000100000",
      "11000110000",
      "11001000010",
      "11001100010",
      "11010000010",
      "11010100010",
      "11011000000",
      "11011010000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000",
      "00000000000");

   signal ra: std_logic_vector(6 downto 0);

begin
   process(clk)
   begin
      if (clk = '1' and clk'event) then
         ra <= a;
      end if;
   end process;

   d <= rom(to_integer(unsigned(ra)));
   c <= "0110111";
end arch;
